��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�
TB�(+�
mQCJXk�ɒ���S�H��U�(�c�H�u���\��֔�PW3�-Ƌ�!���A{���X:��fu��6}�#�����X��/IPz3���y�.w�>u��6�C�
8�x��^.Tq����rF덷�a2vBv���!.d83�,��W	r�����w�NS�kYM����l�L��}�9	k��<�>R�a^e�&�:�*�˻C��ᮮ��n���,��B��m�Ki�1������+�9�D_A�=�1�C�Ͷ:�8�:?����#�M�(�<V]lU����%z��FoTN~�~!_�`%��V^�}�����u��q"��*˫�UHm �uz�Ә����bKr�]�6`"!j�Mr�����Ī:]9�X�P�UJ�����(�%���k��!�������YSJ�s�ߍ�k�J{�=�Z�֐�L�"7�P�� bL^[�J�����+#_9�S�j�QF��8��Cqe�b�F�uVtjC�N�� �K�AC1�M��/R�mψ���3�e�GC���J���Um����(�i���Q�gcW��e� �1��Յ�y)��$+ ?�'�'���CZ��	4�2N�v�@�$�䯕{��d�QP�'A�I��}��{�_��D��+�jɪR&��>�#Q)�5�b?�,�f|��__��
�o�x$s��)�l�w���gA�S��F�X̖�B �Z��e�,̶q���b��șdM�E���V����`����h�~�:���a� �dK��&xo��@'5 S� ��������h�#��1ί��y5��9��xG�$|�m:S6iY)��3iE�^��4�.AɯH�g�ak�PV�~�t�ѐ<������:OC}au	��&z����<�|3o
�(��s�	��{A��o��s[�-,8g�:�ڿo,���5���X_�vWof�,47��y\*W؆�LL1��mJ���%��X�)Q4���fA�ʵ�|)Q=e�L�#|��9$��6^;�N�=�d~��: 7�n�'���������`:[\�H<J>-G���Y:�;�Mri}dq�5��/�Ḝ�T`��^���"?��{�8���%��$��=�f�fV� !����X��
˭gG*jBMb	�������z�f��o������$dP�sL�ڐxn�ڶ�o��.��a�N���|�dҠ����L��<�bnU"I������4o�	�^H�ԯYFDYH�W"��A������B�W��6Ŏ� ���.K��.6��%*Z�([��0�

I-�-��tg)C=D�K��5�Gd_Z�B�=zN��A�J�=7w2�}	h�͐�Gk�%eh���	)Q�$�Xw�h�S���ǌN�61����ó��3�Z����>�clr�O�*����
�j>T?���LB�Y^h���;WMWӀ̈�n��]�piN ��q[�J���z�Y�}CoG62"�x��0`�\8�"�ӫ�cmN��#U^��;�S���!I�aÛ���^̙�v��'
�1��}�{�3A�
�������1��3��{��J���k.'J�*jP����$��'�[sQ��3�1l���R1��v}�F���U!�js�#f]�1���Ja۷s��̊M-�@i�_�^���]T1@�J�fҬs�G��nZ���\�
r� ��؀ߺ�kk�^�����UE�NM��m��yL�=����-��"/x����n*3� �@7Y���b�N�X��ܱ+Cqg��n�v7]���18�듉��P?��t��W���	qJ�}�=��+��Ia,��r�^�]���m�y��;/H��{�"x�s��͠������6\�J�I�D���l�k\7�.fBÕ{&.��
�JB�7f��-��Y~��,+�i-��~����&�~��G�Y��:�O�5���D�N%����{�n�n5��^�	��>w���I������:r!-Ϝ���5+G��b��0���[�^{A0��h��;��&�ਠ+Z�0s���{���Hva�oI=��7��l�D�X�	�^�%s��[�t!�Z�f�(�>��,����ܾx����H��m��>a�� �U�F��U�K!�>��^1L1\@ջWE�nc�Z�I��j�<�8�����?*�����v�'��:�����.<�HV_�S���*��_+S�H�/
��])e�)�Ro y�P�2Æ��Cq���(��1?�DC�Z�3q񐝵��XNϙ�L���=�j���M��P�Bg�|�9��8�9W�/{. �c�-%I��ORG�</Hvh�� �;K���/	���v�{d�wC=t�vo}�D��dIG�~���iل�� #�d�Е�����_:�g,1�	Ϛ�����u���9��K,���\���Մ#�?φ&��W�͌^������2��Q;�䠴x�اJ�u��CU�����:��8֤@�^�O��(X��p0\�j�0�چͽ=o�G���<a����Ui
�|���+˒��y��G�Bx�����oa��v�>q:D��Q�)ˤ�(Z��{���y=�j�;;�R2A"��}E9��hS��S(&G�AM�؅N�^��5/��ɮь`��n�����`q�M�T6��L�VUR8��ʽ?/�-
�}mv�^�����g�	����i�ϳ��JmTL��F�e��m�c-�
�&������sr�WܓҘ�e����?>~*r?�R�LG&+lW�&�N���i
C�p��y`G�om�����M4�G��	��}��UL�I�/I捈Ĉxz0�%a��xm�^|0�����G���ΣP�ͤ���.w��ڶ�;{Y�MY+L=E��.�7L�㣨��W!ek�JO�u@hR!�I�ƁR�Y�z���Ρ���d��\�^�S�:�6�6����N|���rF�o�9s���?��d�bc��hV�JO�IoS�7����J�Q��]��wJ'�S~���|T�xȨ"��-�l��U�3 4�>��k8=x��

�+�N,�+g�9>*8I��Lr-�"��!�Jv&	��	�@$��48Qj�k_���qϩ>ͽA9�R����k�@�i�~�;����H��1��4�mktp���� K�L:Z�F��`�Ew��>8�(��Z������mn�[�m�{�י�O���;.Pߘl-V<
e�r#�7��AI�;�>����.�ӑ��n��K��:j�l��z`�-�M�O�X-��R�$���>J�em@�M���?�+H�#�5�����rPۖ&�i������� ��K���*�1�p �P��ay#�+t�ʔ��~��d�~��v�<H��h�e#�L'������$���c�z�S���5#F�u9תِ�o���8�i�~4�
T�fV��;���?��E �����)�"�*���O�s��!�"]hoS���!�uz��b���F�$�^��c��}1��A��(w��j2����[I��7Nw����5L���q����Ͽng�\8��dJG�� �<5�E���*N[����ߩq>E4�F61K6!�R��.�U��6�?"ܝ�^NІ��(��0*���^}.�Gg2��ԿC�����'H*���2�|���4|�����쇚�е'�S�aZ&_���-T>c�6�t>�`^�r�$>Q������_b�����0��h7��shI<EJL)�AS��a��@fR]t�3�g}S5�,BCf��W�8��[.�c�ZX������a
F������E��q�����޺<�'�"����CY�0G#.�9%�(�%��J?��;��OG��z�F�H�3��\��ꘫV.��� �k;�$��u�p�����������_�_Q��C��Ӝ|:���\�k�*d����<��y����Xa��B,�*\Am�$�;,�=�T�|�U�V\���.�r*����"k�Pע�5��XQ�?<�^0��� �VIn$`��IT׍��V���[� qO|�sa��[��a:��d#�1雖�n��&�W��+��Q��*+�А	��㍧��nSr�ׁI��A �x���<V���~��T��t/����
0��48@��̦6�f;��VN\�x;CD��8.�����շG���aИ�Y�ed�����ew,�p?Q~Fځ�)l�X�k����w�e3����v�� EjS�H�-�d~kAu��N&�W�����Т�i�p�]�)?��/�"�苳
!p����-��V)���$��[nS��9�:tV���"մt;�+�j3�5�AԚ��i�0,l/A������\������0�9�2P�vې	 �!���A�kPBP��[0�����?����U�X':�QΘ-n=�L�%>w�5�(�(��߼��:?{I�AO~Z�e��ǿ�)+��%L�v �8J��Rs7��a�{0���T7cp �F�e Zh��8B�f�*�~�����e�͇��V!x���J�ؙ��rUU����1����M�x����zz����܆�+�Ԣ��9�;I��md�Jd��?�_�P��h��.q�.�
5�c�|T�F;b�K�@����v�j��I�_q)������ǟ���0\�.���(V��ǇK���[R7�?�� ��E��]ԤN���r������vR-�Y4@�>��T �s/��og����0���?̔�-7 װ�St�h���ԍNu�]&� ��-kS����x���sE��vz9��/�e�(�]ҼR�R����\zǰ=gi�??D��xIuX%3����GVeW��ZG�I����2eF�K�p����݃�I]c���	RƘ�|ִ+�]�+w_D�>�3Tz��\"1?s��r#��N��E���n��Üp�������}[n��9�w�.^���f�/6h��E"3����f�T������*]{؟����7)���p!9�E����"0��>�a�L����2�3F�+HG1�Ƣ�}���*�w�W�W&W���c��4��Y�F�ڒe%�����On�S,H����Z�ԵF5m����,)V-u���:N5�2�݆`�B�dA��-�̋��P�}���=�,�:��e�!��kv
r�gs�:��QT�g���6����0���N
S�e���ĭ�Uv�b��'I:S�f|��=�9��Vsm0�xf兡!,�:���ɢ$��W�n�����w� ���d�=
���*�0��/B�>vyJ�7^�\���x���� OM���2�dۥB0؍\t/��y��A�;���g
-���g~���P�#@����.F�i��!_ߝ�켵�a�.۝׸�&���H�u V�
�D�k�&�������t���K��Cy4E�ş���Yj��HBR�|X�R�PA(�c������u�_Q-v�k���p��-�g�4
d��b����,eF��%����%:��v,��ʙ�KӔ���v�u|����=�Y*t0�[�1�] ^N���rp;���������L9g��4n���N�^\��Q��^�7ؒ�.B�y5�h!(p�0Ro"TL�[�'���[%�_��� rA�����~PI����:	^����?T�h��E��@�ē$Z��B�+V7�����b�/�KUz��i��_��4��#�������4��ۋz��n�'�X�|<��;U47xK兓�v�N���A��#jꔰs��|��
Q�) J��Q2��XC٥�q�wJeߋ��%��72P��#�������{ ��ݷo�;w�>��7������Q7�]V3��WUiơ��|R�����r�.�r�1�@�k{P�R���_�v�:��G�pq9[�e��+����.'�A�f�į�+�@b?�c=g���%�=��V��2����{Ĭ��e��Z�;�$c�,�]�J��|5�<EAu��� �2�4�e+���n�M4X��%�? �"·��!_���)U�h݅�N��L��)熓��D!��K����.�w?M� /��u��oLa�⨘T�H���#�l��KŽ��h>�b����������ȌD+���j�� �`�oi�j�h�y\�}�>2V����������a��1 {i��?5[<��7���d�)�����à@�b쩓5w.K���up�'�	�" \�Z�⺅���c���wV�C-{��;�b�Tupѹ���]`��t
h,pCGI�i�ʔsE&d')Z���Z�	\�ٙ1C��e��kE��q�w�!��f�mz�U.������28��N$��Ur᣽�sK��c�E=��]z�-�P&*�&��U�&��gi��ߪf;�=P�X�Ӎ���0��͢������(]���}���4~AM,y�ѫ^⸂q����T#CI����O�DƇX�>�LJM&E�/z�5�.ɜ�!��*��2H�����"d�z��4�q�ADiH~��������fP/����!�˛>���Ҽ�2"]��$��}���D5�$W������$	}�B�c׌�x^u-#,���n�S��`���٪m�}+�c�@6�Vlj�漖dƛ{�):PV����r�[����y��s���Z,�k'��"�u0�P��/t�̡�4�0(C�ӝ]k|�v�|�:Q�L�pX<�k��ET��dۥBM�5�����Tys�8�>��M)Оџ��<pN��n�!���
E;�-�ջ����`��l -Tg�S��ߣ/k�����Q>돾WR�7���`��L�6KVv�������_�f����p��5#BT>��+>7���\6�� f/��]g���bq�2���As��=9�o>䠞;��s�~,
U��H��a�i0o�:N�ɼ~���.�P#����S��_��Z;m��Ǜ>��'��Z�+O�mf���H�t� _0z��>�}�I�J�H}뙱(����s��56�e��W���(�nz���fr۴��X�!�aSv�;i
R��qī��>��z�x����,�e��KО
?U͒�QP&�QÛ�:��%@���g	,�{N�^f��8L�`��������~�(X�mZ�e�~w�q��Af!�H�".������JS��
� �BA���N�U�~��X!�L��`͇��4v���_*"ܺ��O!�{P��S�|��D�?�Ef�Wtd����-��5〡�O��O��Hwdr�}�d��u�p�7��ȣ�W�|*��:�̛'�B��-���qp��Rm��[���Ò��>)�I@��c$RW7��%uDn�4*�\�>)�q,���d�s`�	�*�D�kF`�������=�՘�C�s��xY���2A���K#��_��gi�����H�+y�;��}q�P������TV�Su[�a�z�"e1�K�z�\tݳE!��"�{���Ɗ�����I'����e���mD�O/1P��%|�^��&	)�]��ϙ��\OTQ���d�aX�rq��@�Yv��ۗ$�A�ϝ�d��c.r�z/�U� �P�o?W~���	}uwR����v\�a���ځ�i���6�AF� �r��~�Rh�e�eS�&��R��ὠxm�Z]��KS���4(��:��B7�ǚI΀|�x]l�b� �s�%U*�-�&�׺��qpy����+�h'm�;�i�G2�&��G!���(��bS�4�DAǖ�Η�XX�1)8��Tȯ����躒�/Ц��o>���j�Aȸg� ��T���A���(�f�u�Y�h�-!%��PWS�*^2�\EW�eXu_�&Y��\ �!m�V�)H[�P8͜��qS=F�z�V�n�Mi0��y������73�f����@��N�UKQ8N�]t��F��\kG'�j1�AT�j�9���oCf�t3�Q\���L�	�Q|5���Jb�%M-��@� ��#�fc�� 4+D+����׹�u�����teiڣO�G����ćz��l$Q֏��D�t5�y϶��1���f#J]LL`Z�Q��(,(��6D��I'�^E�̯Ǽ��y+󍇰����l4K�V�!y�|���2،r����2tYΟ��FP�	2��b� ��E�ft;�p�R�Ut�v�	ƌ���U�7-i�h#ߎ�3m�����W%_,h̷���!W`S�����lx���ƿ�J��<:��>K�ס������������zL�g��Q�-YqEa�����	X�����pWw[�>L��� �/ǭꘌ�4�Y��}���َ?�>ɕ1��/�C����rH�dS�-Z�g��ܴ�ڥ���F�"7	�ҍB;���S�_q�/����M8	]_ٜ{��B���8�V���4�ѫ��DցGꊀ�.( �OE��o����'r� [����(ň41!ǥ\��)��<)���cH����X!��,�Fr?E]��f�QZ�?��=�:~,�h6��zr�E�ZL4\���h�G�^,|K�09!ڇ.�`(,�n�'�=6�'���Y#�ֽ�����ⲵ�miH�K0-V!����(^��k�z��ph�>T��ҹ�c�@M��g�Q�eR��|Ź���U0!���3c�5���q�����D����jtYb[�RDe��91E���F!�1Od��d'Mϋ����<е=C�du���8�`��/`%U�j�G+��V�
5����u��_�3R#��Ȯ�O�ε,�dvo
aW5^BaB�oů�}L�>�>4��� i�I�����⁊�/?g�[	��7T'ѣ���A���wM�Gu����'���C�E���kMd�G��fە�����_oI	=H�N5��\��@��K��-�?V%;�L�)��Y[�=��<��+��ܣ�/�S<V�X���n��ϧ��։�8f��j��KQ��al�sD9	)W��@��� �����|:�P>�	[2�������[p �q3Š�Ym2_�yh� ��G��N�'���Q�����;ӱf�sƼy޴�h�D���s�:V�	�.���F��.`�8�뇟O�HWF����n�t9?�[�-*^b+���[�ړ*��T���iVѐ���VI:��ʙ(:K��գ�j��`\����T�� [�>Ͼk�����QnF�ww ��]_I�4�C�*�:r:�.�5L�V��6_/����=>��1��.��Xw�9a{����U�')��.���7��a�c�e9�_��ʱ��㨛u�Ŝ+Y��\ˬҾ(6J��� ��^ly�'�СC��x�Z1�^�9ك���k�`�0���{l�N��/��C�-��h��?^�v*��x6���֮�]��6>���::�Rm�ay��}ђj+?
.����@��UԵm��38��>��������u�:A���Z���0Kw;����X,z���"���Ռk�l�����V�E��F�F��@�`��&�r�g�u%�s� i�[���Xg�
.^�r������u�tj"<��*z�����^| �� ��������$ì1?p$��1NǥH����ȣ��T���\���j�+��7�S�<3
*�3:m7�`y5�C�����N�m�W�OnQAx2�Z�P�~�G/��y(�a +��*���E�b��B?���}x���S
l�ֳS0����$�l����Rls�u�Sǆ9ʖr����8?S���3:�F�����_q��aSkb��>9tUPJ
D�x��χ�.nni��G1���kß%���5 �D1V\��5G,�~g5�aoWd	�+n$kѵ�$�gy1���j����G������g����c�`X
'��Z@:�-l��%���Chs�:n�g�C��ݰ�-�p������=_I����3O>�o�j���fl]�瘜�
-h&}�rW�q��B`1̌|����s��j h��͹����|���P��1y�+�c�ت���_ EGך�+��u���x�G�B�ɤF Ϲ���f����>�c�7S_�TP����W�9i�R�*�5��s�n��}����ݶ�2t �S��-n6�,�1:j,<Z�ׁ2ϖܜ����_I��W��I���3TmCk� 1P�q������WB�V2�E��&�F2�ښ�tƁ����&0_�Y���vٹ��L�#�`��1���b�؊w�(�O�٠�g{�c�9FR0�H�]��ۼc#n��cHI��_Jj-+9��^��λOD���"�LY�8���h�˷<2h�����f�L��Ԍ�JmI��:Q��jv�ղ����X�iP�����>����Vf��!���ŗ���9}1q�u�n��;:ʉQ(H�6�R7��jz�rA�ވ�H4(¯��
i(n&Zzy"�H,(���ʺ����HҩN��$Bp*�QM���HY�!�A_�+�DJ9�P�f��?���<��aڊ��ً�F�мS�	���렐��K�SJl�XΛM�V�]?orx]h(��7��?5�2x~<F� �z���:c���=�khd坙OJ-�ozg,�εS	wX�0l|!w�{�b�O��9\H2<@�����������vNu�ݹ�ȑ �Tz�r���w�<Ϊ���Ծ�I���J�D�:" e�!��L[�!�nE߬�J����C�����[e��1ƾ�:���_�!땎�&AϪ�#6�)UZ9��2c���;�Lr�b�@$�.�cx�g�� ����Ft�@3�$�|��'0Wtn�j5�ҁ����`K�P�����ϴ�e�_�P5{����5�aqO1�$��@$�7t�6x�y��CW��i�-��y�D�%K*�@Mn��X�!�vQ0<B9U�,$?W�l|�ń��u�f�s@���"��y�#����{Ӯp�b�����K]��{�����|�IB�R�g�>�Gp��Eg� �{�:�h���f	�{Es�	'x�g���Jn���٫
:���h��e&=m�"A ���w�z ���J:9m�>w[ָ���\���7��ԧѹ��[T�%�M�c*Y'��=Z*`J;  VZi��O -���E����?��y�H`$���I�{����T��4#�J(������d��y�y�dԪ��#�\�=��(R�7��%!�`u�T@܏1�Z�a���A��]"TՕ�k�LBq�>��8��M��͖��D|ŵ�֍���
�|G�2C��2��۹����������KW��o�|A��!pu����J���6��Hvu0F�$:@g��gd.����-Vc޶]�z����p��d�֕�C���jK��t?�0���S�������:<�d��)�ެ�:����"��-��֓��8'�f�� ���� �=xn/�h9�Bg�~�ɘ���,�͍�. ZB4Э��~��V,mߣ�" d�%�N�^7�W�4��K�`Z�4S�t����7\����RL�+bD1zYw��`'�b;X��1m����+��#��������_Ҷ�~ñ�-����؏�7:"��W��,�,������h�vr�^��ճSek]>
��k�Y��il�c�����J�_�1�X�!`)��'��gU�+�V=��ET�9f%)���r��53�1��H�A���5��E�"8�L�h�t`M6��T�0�]�s� K}�� �����#���k�B�#�*Yk�(H�Nv8a��峭��va(se�D�<����f��c���E<DT�c\��F�� ������AĮ��i�d�� �n����Ԑ6�� �p!��aD�w��L$�n�tv��H>i���`��na�����	�S�Qx)HC̀�dyf�F�2^f�Az�X���!+�}����~
5�A�pM���kA0�4E��� 2ak1^s�C���4 �Ѡiʳ���,P����Q��@�:����?l=�zp)��R�T�%5([���a�X|O����>��I�9�����KY� � ����hهc򨥏����O�H�r�.}J��yt�&:�6
��v4A����OC���@
�r��㣻 {�{�oR5�a�a�@~�p	D��$S�Ȏ�z�|ޖ��H_���1g��k2ĩ%��/庖k�bj(��,nkӜ�8�a¥�����+���ͯ���y�`���
!*=�[�U�;p1@]?�����#;�Ic��
2����7B��\C�����gΡ�N�:ۘ��&�za�u��$D?xD~a�!���>/��M`�ݥ��6�t?w*,*C���	�t	�������Y>�������w��Xh�^�Yl]1�]���ԕ u�R�:wzz8
�^��c�2W���ʠ�4�+��S�F��{6}��@���}1�,�?�9h�yz�� �PL�[�@�����#2�K�QN/Ul�����3>�J��+��t�p^�6�*i#4:Y-z�g�<?���l^g���\*b�T.�+Ƀ�#H�Kd�r!4�ة�o��;0��'1�co-<�8Y�S%��~���~V� ��*���)�J(`������7�;�U�{k�(DN�Z:��-�5��FB��ʔ�#R�S�A�0CԱ�-.��Ķ�rφ���0<��'�FF��y,��Ek�zW�_3����!j��I���q�0�\�8}��A1a��P8dH�:ˍ��
�r��
�{�O�Q�e(���[�����S	ao!H���!�cי.9�"Ff�6�,%����>aK���LX���n��7�F>��}�T���6t|���Q2�6p���f2�9�.�D��6`eL��%��B̓�ڞ��v�`���+��{�y=�������򪎐�'|�7��^��������!� ���_��22��r��]rCh���o���F�q�_/\�z�r�|�k&P�E�	�^�����:x���u%�d�J4�k�tR�S0�z 
�",�h��ɢD��/�yhO�>�*�|m���δ�*���Zh��A����˗���X\�/b+׾aI�ҏ�(�v�>R*>
�Vu|L`��k�v�A1��`w#��`Hl�&�q�ue�
�i8k�hͦ���T0�=����ۂ�Cݧ�?�@��b�p�(\۲���_�x���+�����Bm����JN�{��!�.Bl{����v�"��s�=2?����D�	��AQ�ʋ{`�{K5���%S�H���DP
��$�	�ВW��s������F��L�	A ����<b�r�v�I[[��%����e*)��'��2<n�֐8�(�ˋ:_�w2U�l.q?u��L�����?��g4&�o�M�wZ������낛Y��X��7�悤�<�h�Y��BB!զ��QkE��b�F/��H�jz��y������R�(�ǧ���.�V�`Kڵ2,�\`�#�Fhp�FV�_Rmy��O�˓h�����vۑ
Q��EA
�����_�ۿy�!G�2���m!N@�WQ_�S�b�d���c�A��[�jR�S"a_�膌g�T�[s1�nC!~E�\竟^)g��D���RE��}nr��P`{�_q��SH���q �d�4(��Dik�໎`'��s�<�����	���
���5WU/;`��24{h»�z�.u\�P�&�k�2��8 ��C�,dy	��bQ<)�{������'�n��e�"��p�_���-8�By�$���9��Q�x-[��}1�T��mG�mAE�������<m6@iSe�!ב.e�ɆZ�f��W��!p{@�
L���a=�{������5x"���{���P����Ԏ��US����^a���)���!�L������)?.Җ���[�֜?ѧ�H%�S�kdl?"��`7�_��R�y]'�z�V-vj�g�<���km�r �^�1�.M���oB,��g�BU��"%�������*wܘ�wo(���V�(}�:)c����t���nM]�Ӆ@����J�,<k�" �]����G� &�BF!95��8�b_\`�+O�]���䳀yn����������5�}e�ѫ�� �I
b0na�����c�UG�Q����s�&���<IJ@?��0�Zu�X�-�� ��)d��y�C�%��j����$��c5�9�*p��� � �7rq����w�͢�#)]�]��j�L"��w=)i�u��t��xշV���= �E��LA��������y��u�:1��ۆ�U���l@�d������:B�N���)�q_�<�]a�C�o�����9�[ �kLb ��(:D|�%�&ձ�����Q�R����0��/)���\1>����E(����Zy���'��:�����_p��w?���\8�R��h	���.��4�dn{��g|3����G�uL����p,�$|�j`� �%/6d$��f�Lj2�?�6����<�F�İGV���p@��u}񛽈=�;��*O!�p$P�uuΊ�$�c�>{� ��c�X���g7�uF�VlC��>~[�����?�ٞX��B��3$C�9R��5�؞D���*K��d\!�s�Ľ��-�^�]��q䙈*��tO���s"��c� �0z�ӅM<~ �����w�А����[�����*�W���6Z7�уe��)�b��)�/��HXH�����@���Y�@��*�<��w7�k)�ݶ�AS�	*�4Y��8���sꮄ
�����T��'��G�Z4&�S�&p�q���'���3m4wb=A�'9�;�G�HZx^2�IlzX˕_>��V�/ nYFB�f���3���q���"�p�^�O=L�Ԏ�/�Ls�c���f���B.(7��`�S��
:��k͘ps͝�h��y$s��v�D�%"��q��w��Ođ$�	șM�;v����,�>�"o���ؽ�KA���F��$���#3��T]ƻ��%[q��jF<�>_�#�TAEp�L��cui��J�=�2d��(���B�,N�)Ǿ���^8��6Ykg�J�3M�[��$bd��]\.��S�i{ 3��Z��h̸M[��%f|��4���%4]E��h��DB�ZU�ʦ���n��w�'6%��v�3�����v�D��;�?��6\���kO)s����W��6�U�
���ښM0'�������2��_4��o�f�G:w���OP�O�iq���H�5T�3��gw�>�s�f��~р�
��5�u�I�ҋ���IϲT#߁1r���t=��5��U�h���.��Va�n�PG�@x��v(AR�Bl7�?-�r���g�?�-���I�r͹�F���XK'R���~�Kd-?<�щ����AG�D,�D1���P�J��%���]=��Z/��"����Σ�g�5R��=4	'�Hl����c��$���(n��s�Y���F�V������\g96B�HQ%�����)���!�"�/�b�������ܬ����6K�Ԍ�#��x�d�L����[��-�����4uѦ+e�!`�T����'0�I���o09J�BB`�)d*t���`RT��cS��R.�*�2�G��C{_�\��B�~-��n̶ �!TB��<���\��Z�H�L]�um�Pr-��$�ћӟB�����J�lt���}=��M��cN�~�W?�t���&N%�;�3�����rh	�Lˁ�,�ګu9h���RtA��T�>�@����{�JVms��Z����b����o�Ɠ�NR��L����Jn@�̭��'��4���P��w��Ҫ���b�D�����|<���!\j�����1���ɭ#/�Ak �N�]B�w6��d��������D#�l������ӚF��8WMS��2�3!�>��`����1��H�8r?�Md7���+�����.T��.KO�R�9!�*l\�pK�v���� �ڵ"'��QBc�����}��J�w|{3m�#�{�
�c��<J1�L���2V�� ���J͡�;��y��O�^��t���mI(�&�s�0�H2�e^0�L�k�>_+�.A�3�Y~J��Y�[�Ͷ/�*m�`�*�;���5{�;_�:�����-�M�=�ʈVZ�g��"�\��k� 8��sĐ����%A6>�x����YWDQ��Y�T�.�^L�K�@Œ����ߑ+)=�{�$�(M3������x���u>o��z���9۟S5�"Z���d�4�v
:�NN����gI"��
�C.���q��[��j�Ń�7G(s>�7(�0�vw��W'�LX����kWUf��\���`��"�5������}���.��c����~��-��_�Иq��92�D~��du&�o������ �{���"]��]9B66�Z���ʯ��9��;3zԄ��l2KU�"�0�Z�fj�ɨ۴��|@>�Cy������RjP������_3�������Ts��UU䤾j2u�2�c�w�w�7�znj"g�N�}"��C.���֤�DhqqNk8��(�^m^d����
�qXҪ�@���$��o}����ȩ'�Cl����\�R;^�����Z�l��@�BzTi$"�i�^!��6C����F����̿�S߈s�l����h�/�r�M�ߜ-�S���?��uVֺR�h���qp)�q+�t��1�$��B(m����񼯊�:z��c>ą���۬�~������6�@�vޠu5�� YВz2���{qVB��-��^��G���wn����e�0���ҦOh�y>���N�>�8�Li/1�"G.�@����M����xZ��|y1M+�P�xM{!G\�}�&|���o(���\n�4�ur{l��0l����#F����WqЃ)����=E�����˺����y^�T���L�G��pβEǄ�Z9��A�A}؃ ��8%���oCt�i���n���m�'����C���n�J&��N�q�T�V�N��)rD�7t=dhL��fN����L�S4���JI��OV�G����V��Uf6y��bS�F�Z`
3�����w"X��WP��Knֱ�P7�=�)�ӡC"�����T�J����m���SDF�t���7��,�8M�]Ǟ��Arr��W��c����?H+.t&ĕ*�S�ۉe!�-!���~������8���x����m�[&�awi�`_���D @~�"�Z�FѲ����KNR�b�����%h߉�e�t�� �Xsc�r�?$ n8���u�x?8�}n�����{T{�Q���d��:o�Ԡ%�0��Ql�-�b�3���#��'+O�R�|�_n�ˉ�K�Ù�-O);^���E�*٘��5̨��{M�$������Ox�O���)b���M
L������S�?B�\��C���	��>�#���ê��x3����a�S���*r��[��ÂX`��1��t�A9hO�\>�2�19N� �$n18��'��!:A��c��N�}x%��1w����=<�|��7����#]��6Z���ԓ��٨�-���w��Q8Ǒ���M^�^ޱNm��cڤ��\㩦�hE�3C�������S�)Yo��0m��5L��� }V�L��ʙ�6��S��q�4�Կ]G�:Ff���x�0`5��Mn<�����ڠ(}'�p!�.�-��(�o����0�<�*P^�+�K��t2�2�J�d_��A����F�����l<zC��I������|)u�a+Uc?��&�r~�J���4_��+`���D�\�R���nR��x��8�W����L����S~
��xk��j������v-W�0��@w��+$S�EO���fGK��,�
���u �y�����T�{a���p����0�O�Y�L��f�nt?L��Ll#wj���#p�2��wU<!������ۼ:��ϋj ��~X�Sb��QTH?���\���o����PV���pK�s���p)_�w��_���H��w��ͧ�P&�����bT�?7h��F̆Z/}س�x�fU�j�����E�T�� %?:G`��?�"Z��n5��,��3vo��^��~o�=����Jp/d �=���{K�.ǥ`�x�	�;09�8�!��<���-���Ti��Ǳ��{�T�;R,1�l�I��`Z}�e�0�=�ߔF
�,i���[�]��t��ϙC.��P�y��%����8�C,��J`��1����w����C�֣R�/��A�@�/���1
2���D���[[�z�K�q������ g�5�ާ�J�Mb�WKl�R��� ���	���2�l��,'�_&�.wR;�`eh��g�ǳ����*	���ަ�b���h,{��6�_=!�2K�`%��B3�kS|�[����6�q��jkH�� *��	ƆK�&��g'S��z
��b��,�w'��+�P�X)Xx�P��t��Y��p9�3��(섌����&�.��i.�������Z�X��� �y\v�b��`�Z��7���� B$�KAs�W��,���w����#�ef}m�,Z��21�1�����A�>)�;�T!��;��EW'�į�N�0VL��0�!��U���8SmU/o��L�ܽUZw���ҁ�y'�$��c������Rv_�A��X����7�b�w��	^�@�]Q���FN'"�J�;K::�G�Z�~x��� G��۹dg+jΌ_>b���{Q� 
���'H�F?Vf	>�LO��6�]���ℵd�d�.*B����i�����V�H|�0�X��c���P��WˣM�>��/P��k$|.>�� �	%�|��:P�@h��5�*�#t�IF��i7��E���Jᑡ^�p����#g�ˬo���j�u�o��g΋(ojO�u��ڎc�m�I��/�K����v�?|���?άb9�|P���ף*������n:;�bC
�!��|+>I�!���
�#�B�p�똷>��Ӱ!��$\QO/���ꇈץ�ӊ�����_a(k�f��<�����xh�qD�0�HH���-�n�ʣ�w�&ڈ(SkC�ٍk?K��l��"Q�����l��*�"�� ,�E8���[iz�!%U����c��qT�+<��)Zsn���_���I?k�S��t'|����+K��.=�{�h�>���P�.�S�
I�0׳�"�]�B��H��[UQ�9�
-Q��;��p�����%.��P��@)�X��jgew٫�h�䣦@�7���+�=*�1$lE��GR9F�(�cW�S�M!���W�g�K2������Q���ը )}>X�	��+��:�T��2Pb��4>�����6,�p��c��i �b���1�7g���뵛���f���w:I��z)�J�\��EH��XK��	����ɪ�]Ff'�_�&��sQѫ�'��T��}����B^���jO�^����2nuZgp�1��)�~���3��e��"��-k�PF�q���ڡ��3�^��t�hq���jo�!"ͤ�|����\���?9tJ&e�O�XK�&��:�X�N��㋝������JN�oV��Ϙ54�pj�.#\,��`���rϖ1}�,1�#62EŲ�>o��0�a��Z)�o��^��E!���(y��G�<��(���2��ˍ�|��@4C������X��L�v��m�6M�n������-�dh,��P��$�5�TPƩ!|T�07^=�޷n/�1�샓c�o�&��zo�������U6�[l���1�֕I�|�����f�)+�5�gî#*S��ͼ9��C��y\��=U~MG�~������p�=BK"|,S��<�:60L6�kf�ow��)��:�$���ѹ���˰����]u��7v:<b����U����Y��R:g�����b�q�(�r�k� �c��^�`t~@�ݓ�!��h���JU׈�`�u����?4Q�Z��쓤ի%V�%��=G���
�5�"�3DVЁս;����a�.�~@������V�8N�)[�ooᎩ�Ik�o~%'��3�>�@�ĝ���bY�=��G�,�
�pH4�"K�U]�������#��k7�T]�0�x�u���]���5�O?��5�j>��W�n�ؑ<CO�uA�h��F�k}AI]�jA>�o>�����c'0�;�C�[���H#�ٱu�b�,J��b��{#}p��Dgt�x������.95�}�6?���9w�ͫ�˦�h!~�6�ᨚ��Y��{�����^��M)В�As�Ν�^��ðׂ�Y��^��}����V�Hw�I
�a} '�LCq>*�����u'��P�\�1z�1|�=��ӥ �P�:�o�q���>c�X\6�|�� �%f����^RP�6g8
°2���+���n�>�����F�]�A��Yy���%�ma�K>��>�����=�	�c�Ġ�D{�;-��Pyt^?�`d1�Sp�:��9 ����9��a�3�ô��q=+E��f��l���0F�T{�z�/��N����Fs���栿|��ղl���@$O;L�h���[����lp��5�E2p���؁ �����nRV����H��GG�I�1��3�����!*t���z�ch>���#@����׫�u��g�����LE���S6�|�i'��+^}��JR2�K`�i��|'��1� -��7��_#Od�ST>kSm �G� �
�e9�<!�DV,/N�4��=k�H��8�"ɻ������qc��!�/��S�LҐ��R��G�v����5��]6y���э�I�]��;I��������W4� �o]����N�,��B�:&��r2�3ˣ}>��H��k��a��'Ԡ'�wRizq���h0@��5��G�qun�x�)��G�"��z�?Q��p��^MCP���@�N�$����`U�X�o
�xV]��͹"u�K����a����qۇk���A]S��#v������}P��鲏9}P
�{�*�E3-�������%�9H�{�zKg��N��}l
uX�G��D��v���à��n%wkI�HU;e1PA38D�BC~�΁��h�R�}f��EJ����>m��yʒ�ǰ�9��瞮Cyk�:���p�X�gY�u�T�P�"�[������	-ف����Η&ڞ�
o�eQX�	�{��?\Z�(��Z��Ј���l5�^\��vI�x����祼ưK�Hf��$������@*k<@.�~�[����^�/)ڛ�p*����N�Wk�<q�P|"�u�͉b\���zQ��2۝���:�6�^8��3.�@b���=c���.��ePs�?��P/�`�^L-b+��Vm ��=W&���є,4|�&��n:���MR���z:	�����bi�-�Go屷�wf��[�<Ǽ2Ԡ�����)����M���! ��2�К�c�K��*��P6d���i��ò�Z&��`��c{{��V����v�x~�1�X�����㓛�^Wz��tV�c��+�F�����bT7�v�+� ��6�d��Z��?#�4&����eG�D�3[��Y�3;��C�V�+�9�+ 0U�b�������;;8�!9����޽-+�y�1O�ș#6����X����DGn���L���A�+]a	k��s��IV���3v�= �R�;Ǧ�<x`�/A��H�C���ZT>��Q5q����U��v@�x>*v�z���4Y/�$cnw��W.�;�Qf�����7Y.P�3�+)����:��9˲��a��)��ש���	[?)W=8�h
$��B�=� T'6�	g�$��kJ�ɝ��
((���%&�{c\>@}	��o�G�����&�T�ADà�{�0�����@L*�e@��t��߅��R� ��U�
<������D@'��d�F�2̊���6��b�j�[�g �a��
C���x�/�:*I�O_c�/!�s�� kl>��TfO�4ZG�Љ���	sβ�!i��q�1j��y��E�l�3T� :�����x�>Ϗ7�C�Gf���区z�go#n��Y��X������2ˌ���N��%��ٞ�!�5hX�)q+�;u-[<�b(A���DAsף��po;i����=cV��.�GW�{1r��AĆ�W�A��)\��1`��J�����R�YG�<�d�3��ls�p�N'�Ok�8Pb���(�`�$�N%�Z����"��!FZU?�lX�jwF�5x�)E�$!�3��J��
��Az@*�8���35Ni�֛�@7e¹P �Zs�b�8%+���N�b;��-\�wL����S#\�g#m��|��Í�'j|����+�c㋎�n)<�q���}���^d�K�'����>L���2���z�|��.ʖ�2��Stgk�� 1Q����8uoߴ%�{���̊�k��f ���+[�G�h�nZ)��۠p���>G����W͒yESǌ�Iu$����l���-��-��Q;d��%��9�U8�6�ɣ!Z'UZ�=/��g:���ާ?��K��\�:����4��S*&�!���Y~���E�U	��q�~�����`��as&����Z�/^ʭ��OO�]�gI�4
����}��F4k�i�(T���`PPԬ�ˉ��V���*<�T3+f�?�j�ɍY�]A[h˖�v0�����s�k��LO��u}�<(��N�	@*�ć�*R�
�ՠ�W�����ޮ,��I�������	�A�J�FQ�S����D-M��C�#e;��f�T7������{�V4��z)GR�gI��p��i�xLT�v�lj���2�(W}�TqtX�sy��vJf*L�F+��GIa<�c�e�o�%Z�ѷ`C,Z=�`�8��E�q����y��5�l���_C�?��m�"Dj�,�x�кb1���Ǐ��y�a3O�Pܫ�I8��6�Z�!����v߅��^�M�{F
�u��?�����6e�׾{W8+�9	qD�u�~ܦ#�+�d���=ol��9���H�>�ow_C�~�cU6�	J&`�;b��.侎�ф3g�M�Ri[����]�f�+�OB�Z�#���\T{��fֶ��P>H��8^��ِC;C\O�w爉܄��A�/ȵ�����K�V"���0��/�靌�88g�c��'pgZ��� ��'�k�]v�^{���ax��gq�y�.�^8n�=��՗�Q�n�OqU����t�T�P!?�H֐�wv���*r�� �P&���� ϥ�ER��l��~�_��|��o�^qOa�"BB��xW�G���Lؘ㸃���> G��d��S�O�.�u/�P�H������=�C���U���{�>��SA��˿"��C���VT��S�[J�=ґ�E�=��1$,�M%�����W�Z��%��h���
R���U7|��|'�k�2�<xleD+�ȼ[1T�N��w���G���,�Q[��L]�dN[�P� ��ŤU�9���YJ�u��W?�������^���̠1��c&�cPf���o���"� �� �ʋW
4%��]RW(������<�9���; f��q�PJ�J!HE)/5s��wE��f�,��f�oQ[ r\au��'�y��a9󖁝�5f���XM,���Jb�E���Ȍs�e�ё�W�kυBϲ(;��-�Z�&_Ÿ�3ہ����,0��8֣4��M/I��HR��a�}��cl3��Je��M��W��.k�G���u�5���3���<�k�R�����ҷa?�牭7�8��@=�n:��0Uj���
�4��M�[�R������kW�E��x-���ɞ�yԞ�Oj{F�ۨ\ٔL[+��'!'|�^�
� <5d%�3�Y�'�O!�¸D^��-�~/���L�j�3W�1An��d@��8��/�y��'���K.|��w^�������[���)@D�aqU����!��L�Rx!�'|'��iۡ�Ca�`RV*	�V�����t|5���S{g2�$��^�r������Iv+D������޴k��	�\\�Ϗ�Ө�16/k�@����]#�l�J�I��]�a���(�&�{�(��/^�]�E��i��D#��r3A�w��8j����,��M��6�����O����)h�Q#Dc�9#It{qo��`�0V��[k��-@ ��n��7�:,�R��`4w����MJ��IR�
�>ԛ�q`>�IsPa�XZK���b2�K�
�����^��:�*A�;�j���̢M�;h^����+��w��}��Z�90U����h���%��ۢz�vE���o�<ݽ
�D Y������py�F��ڂ�Qِ�M>j��
4��	�aaL��2�7��0�'ʕH�.��xv0[�Ȃ�ň!� >����uc�&;j}�/V�YhG-���#���]�OfG���q��v'up����?(�������wT
]�j��J����kXZ�*���2�0���ΣF޴�_e� 倩aNY��Ka
ӡ����^�u��q�#꿣%�%A����9'%F`��Fo��^k'�m���5cEM2���W�_�����@9e��f$��J��Ԏ�㦪��J�KEሸ���}!^����q'��þ�h�M���+:kyȿXﰞ���qV����lP*˥!��[��c�uz�[y�48�)���T:K'1x���?�����KËk�9�q��b�ҋ���j��ݢ �}P�b<�=z�م0~t������p�d��I�FwКq7��:�vm��i#��o��{��('V�ؑ~2�s\z�zj�s�E�Y�ïPۻ�=w\��M���׽�n�Qk��\/^� Ir<��G�l��~��>�-AD\I?d�M]�n����r���y�qp��uhHp��x�M��0B$�_B��$m�g�8�"!,�,Oo��Ǿ�� c��`3n��ڳ �_y��Y)q�ޯm%h�[�Z�ԉ4���&�����j<B�,-Z����eG�l��JF�,��#<����P�W����ui�<	�MP�#vc ��&��>|a��E���g�a�L;�] 0 w`N	K_�"2L��/��i��A�gI��n�ȹS�%I{<R�Ҥk�&�o�9b5[:~����X�@��,ρ?�k� �r��ұpȜa���(jϽ���Y��e~I�&�J�S�����*C{]�֍utu���<���8gM�dD[�{pgѥ�@b�2�3�@gכ��}�cZ�B6�~�qG��ԯ{�=��W��_Aǝ��x[-jU)��w�q���E7�w�[�}�Bl�F���Ւ��=P���K)���[������o��ٷ��"��t[��eO��4�0��ؚi:Ws��M�|����A;J���U����vR23�UVFX��e�����a��%"-��Jx.U�o�I8�1�,��?F��U�c �1��k�3�<Ͼ�c�qg��wm���9!_��.��{G-�I��^�ىn���K�j���7� ٛ�S����1�ehˤ�/�ۀ�O���y|_��7�E\�D��L�����D��;�X��`���R�:Xv�܀��a_��D*���"ڴ���=S�0�JJ#_<�b��_/�:wu6����(qʏ/�r�������L2�iD2�2�8�d��]Dl�M��#��w�t�0�v�f-�|Za`�����h0�rzF.��L�2�x~Ϸ/w_�����Yl�j8�{�]�4ѻ�7�ZX�ؖ&?���1H{h����i�?=�T������	n�_�.�jT>�c�M3���l�xo�|�=6�o��O1�rt4�k�;�\�G��PV]�㘷c����-�r���z8BO�|L>�n����+�[]���&���̯)���ܼ8��k���6������L����3��>~h���
�3$������spߣu��2%�n�R[Ho��z��GN��d ��]�-��P�"�L�Ч �Q�i������ ��ྦ�������u��?
��$Rew��~p��.ZޘvM�:��kL�G��J9<�@I5x�Z�����jh�OCzJ���@���/��}ge�ZO�4b�xG���vE�DD.n�<��P,�c�*IH��{ �����o��iA|���B&@0��Mu�@���⧿]��;�*{*� 	�2ցS�J��̷��"t��da�M�|����hv�r3Mn37�a��B)�Γ6��uUg���Pއt[!���7Y56o!�ƹ��J����T��r�.�?^��0��҂T�@�u�0$�E�1ki:��W+��L��j*�z��"<^��q�.� ��v��><�� ���M�@���u�;/�TH�F����� �>�M\���X���#���I5vvFX�f�:fBF�ϼXy�7X�N?@=���_�}Q��r}��/=cL���>�\}B�F6z�j�x�ѓ�]
zs&�t��|��o�Y�9���ݳO�&�5)���2���>>�h���;p���K��Y(���N��7^Oޟ�_b.8������ˣ]��t�y�b��\'V:��g�����Y�������ڇ�T� @�kuʈ��]fH�9��������WR�Z蚉����W�s��� ���=J�V7��t���n�[s.D��CԈr����W�h����0︣�=s��ׯ���V������w	V�5�;-9'�`7O�iix���Y��!6)��(H&E�θ̲).k#m��.�Z�)3��Y��?+�!��Nr�eKP�-�{T�f$�\Ⱦi�z%��*"=9���"�^�]5W6��j�jj�vԹv���w�NZlyi#8P@�=&9|��&��J��������9~U�������M��:�
�m�İ�͂�"}�fc)�x>S�W�U�%�!�f�qU����~��	�[ v[n�������Z�2x��h�#p��h��|S�Bs�!��H��+%�S�ЎתM�rd��)Ly�L�� �G�?'�	��������q%�7�fc|�%���"0�/z���󻻓��B���n�$z� �)�	g/.>vK$�=D�S��3�E����o�~��0S�p	�۬�`����3�,%-+i�I���%��MK�{{3��h�x^ZA3��
�[)�7-��FD|��q}&m��"h?��-Z�+���)y��#������i����I�+�歖��'"�/~�iv�m5G�W��� ��� ��&V�(�љ�j�^�����ߧ{����h�ǽ�d��s����x3�Q�����[��~�hn���F�$S�Q���g%:�ŇgĢ��='��)x�\��Œ�_�U���퐱"2�'��GK�[
�ا~�hOB�:Xh�X��H���Y�����(΢�?�H�V5�V�K�r-�'M�{>&m��Ⱥ��
��2��_�������]����'tPT�J��(l�B�Fo?�8WJ����/�q���6����GR��f)�C��0F�F�BF�ɪ�i��KL�[/:�}����'T0�A�uH�Hա֦�iq! !6�ջ|��;~���1�= +p�Dnۤ�[�_�Acd=�k��oJŻ�=����!w�UW�Y
�Z�ԝ!sg�2��0��18g�3:]��cAWQݗ�:�T:�C�4���b����Wd�:�GER0X�w�+�xZJ�%;�55!/�Iz���w�}Aqܤ������r�Dw�wa�-6��?��ǈ]e�!䈒%�і����Kjkn��mz*���o�f ��g��߼U�(��wu�tS7gjm6)�_�}>�e�	��CY.�ͩ���Ie�t@��ԛ��"}2���*A��i�;;f���I���������#���y�I�%Ιڭ�v�<�7x=����3�� @5�d��$ �����4~6��%o���f��ˀ�d�f�dS��m?��5
�4���.6A�� N��� �&R:�k��`s�M����R��]}ۇ�W"S�v����g��|۟��ĹzF~fPG��Uzt������<���c8����5��\^��]��Lʚ~m�Es�X���ˠ3�{�����@���Phٛ����z��9}4�`8^c�w{@W&������m7k���tM��+O���@6~
R�䊚b~���,:�ӹ4#zHEjB��2�J�[���y-J�]o��|��)Ɇ��{���A*2|4Ʈ��m��2�?qoHZ(�C[X��MS�[*y'�;��'����X����{��Oj}*���?�mW��ލ4��/Rɐ$Mߙ�8q�C�ًdk�7X_ꓲRS���K�:�UKo�#�\z������]EN��n���n3,h�,5F�L�bv<�b��c�6�${ ����r/E�I�`�{!�V�I�Ic�"�ǁ��-��<W2�%ml �Ey�x	}&Q�d,E�g�����\�]�k�ƛ��\����M ʍ'�Ξ���8��ly%�C��pkf�H(�1�.%j�j����,���\�*����R��fJXD����#�+�}�*B7��c���ȉ���-.� g�B#�_�k�ݼ����C.��)c�R$��Mq)D�I�k[�m���?/՚���ERC�m�0w��iM����T�/�v5
����EJ��훫�^��F�(��5#��/�^w0�!�MI�caHo=$!��	���U3m�+�����thi���aܱ1��ԕ/3��ݜ��IJ���r��TC�b����nOPq��:�fCi�#-�f��y9�����a�s��-Xy)ԩ-��.z�r����"���Z��'V���N��(�G�/e�w�~� ,Dlx�.M��]V*@�^�{����aȐ���(��B9�[>qQ�qQ-���.H�J:�N6vԹ�;xud]���?E�E~�%�|�[Ű����S0 H�d8^q���j؍�=��8�}T6��oO�"&��`��c`��Y6qE������ӻ��,�-HĴ1熭3i�1��<םҳ���:�A�Z������7L������/������f���Ƕ��-�T��q�*6,��DU��T�ݨ�Di,ȱ��85x�����*�*F���ѱ#��f�+�*E�4X����?̉W��O�hp�(�sN�¤�CiMl�����[�� �g�/�I/���VS8�`�K%Mw�u`|-��Y*�r�����K����xe# E?F��Ye�h�1JDA�>T��Gq��1��z3���c��`?���uQ���/@��_͔�r�fY�_���!��aҌ�'��8�%�JVR&"c,���]�I����
?���������9[ڢ̭�̴��ؽ���ك��"#����3�/?Ռ�&0�Թ�w�;4�@�x��7�K�+��3wMd�VyLu�)�BώBG��i���0Xk>�zQ�q�G�n�+�ߌ�0�E0E6y-i�<�;�<�ºlDy-��0��� �V�`H�2^f��1�}EV����;�'�$���kAC�c�'�_u<�/��9��Ը�<y�V�D%�rs~S����}���U�#��@�YP�cG��rB˜3��|�aŎ�)4i=9�)}?C^!m�Ŗ�c��sIxVhS�@)���`���̳��_�O���N��~��.���]&�r�/0-Q��9q��X],�16��r<N$��=׍a[悎�h�H�N����j��<ѩ��<R�J	e<~�UCs%�y�"'��+S��b���|�?����i�qJ�zy�8P�|��:�D`*
���������1�ԯ&�eNY���z�^�y�I8`V�)ت��Q'�+�s��k�ͦ��W04Z��pG�*���^�de��W������L�4�0j���~	��G8��	n�鋿�B���z^aa����o��T(T�]�;�:��3C�
�r�D��8�3����JO�Q�Mr,���2�2�U����'�o���XV�/��'�Z�G��?��a�W��I[%�c�i��i�:�d3�&�Cn�R���x�;�8��[����*FE��=cȩ��b$+0�R�$����OD������ğ���]N-�c֨��z��p6�r�Ā7xC����!ċ��>�&9-��>�S�T��\>��1��FDn���<���py�scK�z��㏻�CD�r�����"7U���yi�!��)j�ұ��q�;?�����2OrM�-���K��V��U%����}Hw��Cr�����)�A�]^�F8Z0�i=A��?��{]%@��,<L��9|z8�J@p~�)��ccq��� uL��!�����8$�ԡ}V��$��K��{UvlcT�Çh��ëu�I�����F�p���@kA�j��t_4u�?c��)���ӛ��4�E����-h�M2b}YA�R����_H���D��8�%�ni½d�Ȉ�$�"CxX;_��uP�3	p�Wv��~�騹F�P�FF��3ۘ���Y�{~ʉ�.�ĭCe{�W��,��:~���V�/yC��#�gN�(\<�Ta��R�'�}i�"iH����<�lq�7�C�`y;`c�/�ZF��6�Q����Z@�l���$��;�l�Y���Ӧ��'��J�%��N���>R"�s����\��ᾫ�
CB�y��d���V��aɌܠD� 1J��\��F�p�pԨnQu���e+�ݭe����tZ�y��J�l�������g�@`x2��Dk-�5Q�!0NPO�^�)^��1������������4!����Q����fؐ��Ij&�Z0p(:�t�Q�S*Я��d�7�?�-'���>�L"�!/[��T����'.�#F|���4,��B]��)=��'Q88�#L���T�Ė�CMe���n�q�k�G�����B~P�`���{v~����Vs��E|S� ����k��j+&(��]�ͺlg��Z��<��b�C�>��R;�l�{��김�yy�,�jT� srkV�G������<����A�ݭ����G�]���W��#Ek ��+����i�%p0ZŦ��ja^���g����:sQ<��ȘhH�%� �Y�H���[�,+(�;|W6�ۦ�Uo�&�=iW_��D�EI��2j-������F:".��Ni`6�����?�s,}�ɷa���b��"�J8��V�'Q�~���B�{#L@g4�k��N���~�gc<nɩ� �?B7��i/�01WY��j2�0�.3�l�/��X���1����c̭����"�+=��\,G� ]�E7��k�.���ğ��Dm�h�8Z��.J"�"xb��9�	���/$�W!͗�p-�\���l���i3v��yO�A�ςz�9��$ڌX���^��*�`�k7z�]6s/L�r�X����P����F�Mą���b4Ζ��%ʞ{'�珸Iw6PE?��s�$F��|�x���,YXCW{\qLy����A�pźG7�J�
���!(�N�l�J��V�|x�~3v�9{B�ԙ|��� ��pH����wbz������=ʜ�9��}�J_a���m�ڳ�8��[� ِ/
�	 �w��sBs�`��=//����.8t�n�=߅�Ө�^��S��L�[�t���kq�I'�����;Yε&II��q^���a��QL��FZS�͇çfTu�w��ξ8�n���ֺ���!;��6��_6���@���d`�Wr0B���=.	t �4�>ǌBK�2�DR���j�"�Q��KVL�T����@��?hPeK�h����\��1t -]
D���0�A��� Fw��1-1�D���3��X������ɰ��#��p���}by��,�F�tR0%��9-Q�?�#�֔�y�P�8��s]�� &fV)-�sˤ�I,(��ME~\���c������T�_�4��ۻ�}Z�I9�+pS���eT����MW��0�#�����?-�q-��=Q��@C�c���P��{ӌ�k��� �8�ɞS2���qF��pF�МZ[���IF��H�[ވ�]��f��e�l�ͱ�\�����fpT�X�>\tOt�W�vy�oa�~��qVz� ��.�t�Y������E������x!^��o��n|
��sv&�A��yy��Jr�Y�'���\���$m���D�$�F�_�f� ?�ɏT�i�����L=l�]����*�8������"���Y�(�����i���Q+�����*�ߡ��&��8낏@u�7Ɲ��y��y���!�~J�������\JWvZ8�X�Qz�yv�?&�W��s0K؛�2�0d=�tFBGw�X�L�m{��no|��.o��!�$f;��fQ����Ä��1���д��|�c�f]R(�����ƫ;�����i)�#ňgNGfؚw�M��(~��$
���F��X��
CBa�|MBVѳ�co2�5dkݣ�)�8^�)�d��2��Z1��<k<���s�k�uo�V�������Y��{:�=^�6�r�o�2�3���h'�̽�͓_�§n�b8��N���;"��"�PL☠�.��}`��C�z�N����>�k�	t���/�������)�JJE��$��ϩ���+Ƌ2�.��� ���J����v�g�N���Gpq�uυ^k�ٿ��0f;̦j�ÄF�QRhO]��>�G4!
�5Ԯ���v�vK�:�$?.aD�5cbN��O�"�y�v0��FvͰ�-ӭ�NNV�D�'������!(�Z����A�����_�f�$�m��k_�#l��,}���i�'cW�BJ����}����Sڞ3�BP��ƻ������i��V?e�?+_n���dHU��"0�g�4�9a�T�H�V?��H�H��aw�ţ�WT|��񒾚���R��hYpJ�s�P0**-:��dh ���V���W���1�f�j���O2A%`ɷk1'2��aj=��MrK�l�8w�3m�# 4�c��#[���L_��A��Uф��'��:��c�16�g����жYq��ʀ���~�^��E�����#�H�ș��na�!�T�|?B8�:�i�' y"��%�;q�a*�U���3�Rt�K�7��j_U�
r��Xii-jb~Y�o�=�>{@vi�{�)e-m��@a&�1��Ak��FqC<�.�_�I���+�'}��@ٝۺ�/;>�d, ���
j��0���^i��@��"O�C�#:tK�S#$ĸ�_q���v���H����ފ��n������P놾��C\I^t7�D��]�'W��'�F�!�.A�ā
�X1�_�P�gA{�P������@���M����(3DAF�4��1��?1?���}�ӊ��0�]�E30��?!�� FӃ�p�� 0�sE��)E�����'I�*}1!U"\���� 땒̌K�z樳��,9����~���c�#M�L�aQ�<۔��ʏ����W.0V�i��Ӈ�߽�����i+^�Py:T��ʃ�;�#=f@ןbu̮�� �t���ƄG�ɜҨO�vϔCz�=����1���U��S��yJ%w����G��7��%!Y)I�E��6��p��4gL�OBX��8�&w�U焃i͂��ѧ�}�	�}d&'0m��U�ӷ�m3{e���/���{/�Ehm�M���h� ��a��U��5��D	 [w�,�ӃZi,Q�BNb.Q��ze�o	���4\ls��זO-D���FV94����~�շ6�i�A�ӱ�3_�jz6�J�������� �9��o	
�T*��[�lu5�:�Q_B�,��Fm��|A�U�
+n֐�^"�}KD��z��פ���%�@t�oe"��,Ӽ`bSR��'<g�h�f��?�Fj~zL2��x�.����W�G����a��׍�#л�-"�(����@���=#��;P����g{p���y{ؐnҐN�~�� ��������n���nD��1_�q��b��C�Bj���;��L�E��e���Z�Tn:��i��Ve»�K�FQ��=���w���:vsOd��Zu��
�4�_x�@WPGHv�X�2�+c��s���c�H���E��=������˦�aG/�	��l}�[���i@9��6zgA\��������<gP��S�����ĥ?� Nb�b�R�,}Jr-���X;�[^[���b&n�� #���ǌ_��Xx�����ghah]�ة!���Y�8|*X�w��"����44�3\Szg�"�67���;��n3�5X�4ϵ����uúڶ�M�N�2�9V3JE s�����/�����RJY�`> _;���h���:��Y��TR9��T.KxY�1�HF�R��i���T^1��q�e�``����<I�5S�Y����p*��P��A`a@~�]�ejV�0[�̌g(�S/Q�����D?V}Ku�@���l�.���k��G�?.t�~G��&l��C��s<�^X+���x���¹e�7o��Ae��V,�,3�Y�e���'�T��nf��?���d隆�LnR�g|d�g�]���D]|@��%��k��-\��8���·�����<���<������O��6���ZowAo$3:�|�Q�p��{����S�3��YF,�V�
d�	�n�TG�3S���Q�"��7P{U̬�~:��]�l�?�F�\���q�B<`�8t�-0ѹ�7;O�KѤ��J!7^.M�0��7������ʭ�1?����.`�����6BG���z����o}0���BOU��lx��a�Uy�x{�at������s �����2c���I��9�;*�儫*ʈ���ϻE�%���%S�xhiT�O��=|k�,� �`XuK,�M�����9��CWz�����˷���)��j�i�1o�i"��|�p#,mo��h OG�ŧu�tB ���\M����︼�:�a�)ҵ� =��;8��,d!F:�v������� =x�r�iK=G���(�u�>���_��tr�{Ȱ�:�*�\ڋ)�7���$�r)Ә�'8������͇�]cK�at��
X����ȄvF�p�l�%$�&���u�GY�$j�%hR)�0�є�U��d�X5�,�'�� ��ޜ��_ͼ=��`�V�
��ǡ�(|`�>
�ʕ%�BA.��a�ʏ��`ɴU��>lEx=�5�����ҕ}�|���o�kex�C���͙
��e��a�x�S�!xv�7�Ĭ�p14����(+�F}/I^s����^�n
����q���4��k�#����vU� {�n&�, r|��1q2*+��t�44�}��[��C����d=�vJL�2Л6�c�n��'0^W�=�L_�H�-����<�'~�d�[DG'�8��.�"<�;���Yo�.n�dQ_�`s�*z���:����<����gޑ�o��oj�J�J���:
*=4�@��D����e�L���'n5~�g����C\k�H.h��j���_��c�:-��_z�L���z�;ʍ�x�:]M�J������zQ>����d��\R�p���ߩ��R4z�Rs�d=�JL�:U��Ч�7��C��~����D�����$���k��vas�Yf$�C��``�Dښ��@�'�/���\ټ�?��$�C��#;�_��h�Š��ֆ�|u���e�>م�� J����4q5�-��xQ�f�#L�B��S��#-�����e���0�զ�adE6��>3j����WSb�(en't�r�i{��[؏���7C���2E�qH.�X	/�t��e��8��я�7;8;*~x>�B�=�F@�dj&��g�+M��9�'!���F��^
`�I��>]ǹ�0m��M��싃NHE;YFf�e|9d�>�Y����$��'-+)k9���K�!�Q���ɫ5:p����F����Y��.�N:���;�@��yx�22Yf>�N	�_�%�s�*�ҵ��X��8�p�Q��Ҥr���1қ`�r�d��W5�.kB�l�
�У�l�@��7Hh�S����s���%M @�E�y"�!չ0gG�l��)�9ܳ�l�9�U��m���Ξ���>NZ�@�������s	h�򮚏���I�����F�i�V�ʉ�d�8I��2�����2r��
�~S�HD��Dm���I����5�K,��j'Dx�%Ж�p�4�Twa3KWvVx�&H�P��B��>P5��c��]�K?�=�_�n@:49���b�@;� a�aJZ�m��0��:=!�3+�<����TC
;����[��|����י��
�G�_�,Ώi�ټ͌2-{�5J�I  ��:���q58����9�h���r���Q}b���,�F�=��-�h:(�\q(!��*\s`l���B%��8F�s:Ɍա��?D3F�'�����n\;���%ȡ������>׋��{B�7u�4]�ohI��j<u����>��A�j�����x,�L5�[YOrGl.v����`ni�[>�fJ2;�P{���گ8�qM}0;v�I '\5�A駋;��.�5�����IB#Qu��dz�	J^��
��Z�J���d0�SZ`%���\(���P� ���l��Nͺ1�xfa��i��T#��;���ip�(:8~���ZR����Kk[�	u+AZ�A� m���,s��5�ECY��H���( ��F�p]�RvP�(��
�$�ZiNKH٩m<훤�;��J��c�3_���;����I�����`�?����7��8�MU�7N��؍0wy�S�3�аs�c{��3Ϙ���O��@��1��t��p�����]�m��7�X�j�r�'��� cSZ P�a!ƹK0l�hR�u�2m36�ꇻ����en�\���<�� ��K���~	��z�\I�W<�0	�f����SPrH����o��c.i\�phI�F��4[�6��é!�L�xN�RJ��s�����]!߳1�S<�d�sb� �Ё����-�8T��qh���Q��_���J�I�P��c�UD��k)�\�~<J�bBE(���XU)vۍ��]H����NY'�j�A���Z)�sd:Z��6Ţl��E�t�^XM7����Q=u�uaX��@��=�
��x.)��M�Z�ܦ�k�칛�&'o�r�W�e�Ft乸��GDG6�Dr�0+G4��9�<�r�X��N䗨e���4�/��{�؏�!<�<�#��K���@�z�K������3%�o�k���kR�ɯ�BJ���y������?:�=Tѓb��A���wO�IB�TZ@����T�����O'��!���xu2�7�A�೫H�D�-�/�����j�����ɶa��ܳ&>��e
����bɳ�
<�N�X|�i�+��ܱکd��	U��JO��Ĕ�����u����*"Q�Τ{�����ƀQ��8[y�O�p�l���w��V({=�� I���h3(�ڎd�l��'Z�
�m�I3	�;�a�N��A����9˴��5lE�\������k�Un�����`�揕ql�5�$GH�0�ʓ��s^���s�\�'��k���˺H�Y|~�?�^�x�����G�Xpn�|L�Њ���D�P�D��%�x�s�stOD�Px��a&��,�SD������"�Z/ (���r:?�9J��c�jrL<���M�>��	Pɚ�ud��Geg9XՀP^�������i�F�}�
�Z��@kYsso2.��K�ƍ�<:�n*$�޳]�J���~C�0�]�J�����H�ƥ��ŕx�NJ��$��O	�D2������21�zqb��
ַ>bYk�+��-X��\�Mg��s�JZ�<��7Z��f�)��$��#ә#\��84׍o����0�N�'�]T�H��^RCm��B���Rt�fCE�B ���)P@@�aM6�h׳F�����`LT���"�Ԭ��)Ly"������]�7�Ӗ�/�|3bh�u梱-q�ڤc�?~$L���{��2�0��%"������ՙB��4�S���N��2��O�?߁�߳����)�^��U�n^ܫ��xB�~�Jk+��%�.�ȤK����C�����o�OLc�6dQFCV7`��+=�FF;9���$�l`��ucX!��N~�`p�O첨o"���\b��3H���6�Iަ��C@
&l[4܇���<�p�����^�j:�|����3r�6 �u�o�D������`��S �h��8��(#r�?���&SC����@I�lNo��81�,�������b�<�oa�dI����=4�P-Wˮ p�����8�H�/p{�̩-r;������$�I�@�Њl�i
���]����a��5�?��%�?���9���$)��Z������!�F��ņn���o����Mew�'1Q#z����V�0n�	y��]a�;���8+�A��vx�0�D�*.+���c��xV]J),H�p��ACr�K��IR�>��!�i]��4ˢ�T#��ɂ̶��	 ��Q4�m�<�k����SQ���}CWzu
7>nnt�I#��]�p,���^h�8N��X3�m��i3c1�jwq��㩌W�Z��X}���j}Gwg��$��u�X�#�����϶�N���sZ%i~g��"H7��ܟ��� �7A�~�M5��x?��5����Y4��;8��qM���w�\��l�X�QbE����$8K����%r	U����񕯹Ǯ/�fF���m�p�������o����H�[c�u�8���4E�j^���6QߚT"Y�02~�;	KQ�㊕��Լ\��\W쳗�є��g�<�'�X�6� 7@2'�����H��y���c����%����]��4h*|�ܚ@�n~܍��g9늠^��tkS9꘻cV���&�n�ښT �9�s�ʵ�:�0)� � �)�i�{ڴ"�Q$��"�A��'����Z�aV�<W�W~���m�̊�"�?aGT=DX��mY�(��Ϗ���ڍ���w�[`몛O�B�C�����F�ߖ������wg%n�:E��j�����+��� ����$�a�`���yV�GCC�a�)	t�i~T��9 �X�s��n �R;Kb\xak�·���I�Qbm����1�
o�Tp��_Gho��D7F�w�o8ݟJ{p���d�p�Z��3~^g$��hh��2��|��hr�^=�r��\wfZf$�@���_4�8ٍR&�_�n,�8�K2ܩ�w5�&�_�6��t_�	�&Nx�"�T)���8�;���=��v@׀����[w}j������x�M�y��tk����"L�t�v�c����j��\#B0��d\kF��GG��ቦx��1�۽f������4�<Jq�K�<Cڕ5�=��R���X��iX]�Dy������2��#G�8l8n���������Q7dF5Zধ�VPm~M�įO!grI:�l�S/��<�.��k6@?;C�{6��x_��E�U��4L���$2`h��W�s�ј#)�����/����FHN$A�{��gO5A��
	Ju[A�$��Q)zߒ���/ԶꃐϤ{�Pw�QB��\�/z�>���ƿ.]�V���0��2��V��5�Dc���ါ�t�������HX���S����FE��\V�ݓl9?0�m�@6W۸&9�&k�F/�|��2�1�w?�W�z�5Е�`!ˮ<=�3���koٚ>CG� ��ɿ�*q��f�ݯ*������E3 ����g*����\}Hgm�8ȸ��T�R�P��[���2�,�$$�&Mt�������2"Y�,�m��:r	�v�^��iMf��/c�Sƣ�q��չ�U�m�\R���0��� 75W2k?>������8��c�����v?:�6�ҔH�)Bj�H��m�l���4�b���Q����cGh�	#MnjO%�#B��}�*>В�l��GO����&�t�7��\�Uu�0� �J8Ŀp�;�;b�����%����)5��~&�z楻�$0ڸ �G�Y:�H2c�����_֣+p��^_�'Z�V�ǂ��8�1��ݶM�����*G?*�6u�"0�*7��%8�3Q�6����{�;dl���`!T&��9��'	��ֿf���}�˞]�YyH�y!B�mmӔ�K(�5D�=-H�6��b_r����H3��|N���(�8����F��8��<g�.��K.H�I��B?��N���i���p����H�Ij��2b����1(��p��l��y�x��W��G�)l�A*��Ue�ӝt(��J�Wr׳�tǠ�C�~�_���+�p蠀ǯs�����^��
>ѽs S4�l�A��v�NEӒ� ��Y�A����m�����I��4q�+0�"�P�>���rG��}��'���tW�� nf��4g�h��%=,0{-f9=jHҺ)�5���G�� �� ��t��x1���n7��D�쮾�\>�%%=z�\��i�	Qk���i���Q�)�O�f��Ն�h/0.cOb!�;Қ�o܀P{�O3x����w�e�z�^X>�;��V��e�~�H�A	=+�
�U���B����M�(i�~2��)��c�m0�#1y��ol���܀�W	��6e�E��)�s�����Ӳ 1
��O��ΠFu^����1^e��ueO�1I7��5e��w5�9 �{�=)�{J��8`Ԭ'}�3��,�8I���76* ٵ  I�K��M[���qj�]-�g	�6�#,8�B��|�9u�|)�8	{��]4[8f�ΈV�=�ی_��$!`nE ) �
���}��a$`u/�ۛ���V@,�ebMU��Q��ۣ�wQ�=�g�c�G���?;�s�G������/�\����k�����S]UHGt��)L�"�)I<h�}����%1�Yލm����0q�g[�P^w�8�ڒK�z�W�����<9�?8���]��*� Vũx/r�osa��fQ��d�⯐�7TdrCU�}�w�Q��x�&�Sh���)�n��G���`�yu[Rku�^��&��Utb�Y�63�����ޔ���o���|�	�F��5Ki�WM�ˑ�Fm�K��k����1W��kQ��i�C��J��s�k�'��5��F�ܖ����'���m��:�I�Ι�i��;N�.��J?{x�/Q�&OLxM��
�����UAN�צ�ƶ,���{�$8���^�KHЦ�a�:���p�m0������v �����%��-C�p��[a�K�za����J"�� ��3�U��[��8�?�B,�B�c���~�a)��u@OՆ۬]��Cu�F�^���tO��_�_����H
!m   �A��+���J�p��7+i���^Xyd�ُ��8u�}V]�qB)��@i������ʫ[��Q@a���	[<-�5�v�)D���Ё���h��-���F��9�q�{�g.�X����@ٗ�7�@��M�� )����D�{�t!�z8���Q��jTò����y^��I��9���jI�� B�&��|]H��^�0�.��[�&��/)�nrU"cH�7BH�� Ar
=Iȝ�9ԲϬQ�B�j���� o������K�/�UdT��0�d��3���E
*�U�juxT����B�pG�ks���,�Ux��*��� a5��#�t��tiI�T���6c�ccS��$��ζ� �VY\+��9�_�6.�j�¿���c6G���^g�ѨP�� x�
���.o������n�Ӊ��O.p�_������y��znG�~Ma�s�Pg\�1��<�/��누�~u�<�u�(�������ğ��������n@�n7+�����"%�
���2J�e)��1ߗ3⽙�P�=i�������&:�U\f6�}����~���:�;�?����H-�����]�ep���:�G#�P��Z����2:R[	0=�G6Cƾ�~�-�U�6�T�]��C9�c�摔B0ͻ��s����*�Ǳd��������.oE��Y�'���(�~��.�_WP�v���^c�o�l�P��� آ��:��T75�:
؂�,
p��3K��ⅺ�w���p�3����}G-�Y_K�qi�t�� 
(�G���s�͗pf#^k���c��)�����l�7P@^ r���� ����E�iDs*��}�'fw�����`+��n��	��$��&�qp�/�C�i��I���_���a@t��m%G_��g� �'�m���0��4����u�v�K�fz?0�R'����vǐ���}ޮ�R��8(6�!�(Z7jea��7��oT-hQG[�L��$��-E8X݄(�)�ɯ�k۹��j/��(yb>#v􌊔C-�v���ǈS-f�;(��T('kWS��.�^/�QS�"'9�l�V��Cl!�w���xf'o`yiMJ�Ώ����xj��V$I+���M�:N�����U��NG��:u��=H�w��i����8�o�z�u�e��p�ދ,��TW׵nc�΋�V�����L�>��Ȓ^g
t�d=�D�e��L���9��wUMi���W�eE
2�����P.��?��U�x8=�x�-���03@��ia�R�({\��k�W��1�Q���fiI�}��`mF�Y`�>��[����"'�.�"��}���^���܀�['8pE�_��r,R����vzB�AIX-��3��c2�s��գ�@;�T�����Z���B=Tz:نm�\��'�I�ܰQ}�Is��}����3`����{��Z�P�dC4�{�-���W+Y��\`-�sZ~�ND�ao�@�f���>���A.Ёo��t��{N�^#qa���p�i*�`�#?�1�<�O�m�r�v0�kIpi8���;@����|�/@`��H���L�όW�ط�ݍ��H�Mz����\��x<�a�&�Ө٤�`K�~G�	��6���|:�*����u����=��b-�K?��B8>������"�W��l�_t�a��6E�T
�FY��X2b�b��=U��7ΉnNyB���_�%{}
Q�;�j6�����Ii濛�g��S3��օ}��奓oZ;.j���6<�Wd1���\2�&DW���4w�G�:��>|"k�;�;�_kmx�8��I�8�g�R��i)6,��w$I����1S4#�x8ًdX�<������@��ٸ�Z���d�ܩ�ۧ���F�l���E�ETfhj�r�*�-;�R�8����l�����'em�E��;���U�m��uGVr�ui�+!W��Z�ܵ��?_G*�����+"�ARCu-���+�j^���g䭤u�*oZ��5JCm�)tt,������JHJYI�,�J�K�A�U�2�'�RE3�U����Cn���p���/HO�f�ə�k���e	�����<���qi�@g31fI:N=ݲ�e�V�h�ySJ5�r���[	�+�P���e�}O.siR�Ζ��F��:�f�nw&&>���_F)I��E���d��hF�b;�5�M�84ʅ'�ڕ5�N_"�0j�r&l�mfUks�o�g�n"�P�x���107���r��fƳD�7�\���!	 5�(���c����,����%.�$����w+�'�C�#�}n���S�2-QB�w�CE��9��
�0���y����뫕-`��ȧF�X ����h����jbt	 K�����! 7��=���9�o�qx���/W'?�"k�6?�{&T8A���X�״�����U*��UKFL�"a$pު:��[4 s�΄6�U#�:�Ү���^�ɻA{��>�R���t�\�)�&�y���_^oD)'.V�,_Bn����q0��H�#3��2�Z0�=�Kx>��C*Pb9-;��5D|�;H�+�5h�Q�AgY�U��+����x+����֮}8����k8��]�|�f�&΁��z(-�~����D�'%V5Ԡ������3Ut����*���YJ��0�5�H��Q��l6f��E�߂�+�
�Qz��õ򍛍�n�n����!�C��9e+�oJ���?����)T���y�J캜#���o�TtB� ����m[ە1�R0g(k��o���<=�HK�3�N����EXJ"�x�43M(���,Qc�;5���W�4�H��˶�~e��ؠA��5��1�g)�ˠx�U�x.�\�ׇ�����˭K��ߤ ������	�w:�5ݿ�ѓ�Z�����FF/�2��k�cn��S\]���QV���%xp'8�`P��R��~���?�V�?_L����1(�E"�+��3����C��q(��]�(q}���p�Q<%�s�����no�]�,ݹ��[}�m\y�bl�N��wf����!=��k��q�`�I��V�X����38�׎fe�^���d�1&A�^fr���13���}��W�/W�R�`
��3���/��Ҟ.�,��l�D묢"k��<L�u�
,�% ��o@�y��!� ���W4�| �����rJ���v������2aϋ~���k�� �(;�&�e��B�t׼\�M���w@��v��t�y#b�n�"�PpH�"���f>�ܝ��4b~%LieG��-`j���i�hi�2"9 ��WEl?�����=�6J��������K��ݨF�~����I� ������J���Xn�$�C�M�8��r�	f#��hI|2W��Z6aⅿ:@��#�N�{�fe- L���h��H��K'�R�_��EyI��դS�"�n8dmo�"D��G���qgW&�fCU�.OI���H<��Ԧ_X���A�r`qgF��7'��ݰ��S�x��q��XV�
řA��^���Q�,��@�ܷ�oO��nm�Xoy�n�ǐ��ԧiw���#���̯ ��
�F�,�Dx6
�@j��{P��'�=�� Dќ�51�
jQU���:�Y.�h���N����tS�P}��B��!���]p��8��na&xD�*Sz��n�>�J��q'�|%U'�8��e6�Xٚ�3G�-{���@^� �%����~�g��Uы�d�\5��G��-�j�ǎ���^��1�_'B�4��Ab rht5�q�nx��`¹� �Z3y��6N��t ����Q���K�C�N��\ƴ���U�|��V�T]j�2��v��b%yA����5��6�-�k]�$y��`WN�����:'�R�!��3��?�^Z�˳C�fj�u��!��EkEǬ[f�c��`
� ��G֪ݶ꽫}<Ó�m��e���-)9�u�G����P0��hQS~&�;��d���(OfI;v�r2�	�S$�nWi ��7_ݰ��`ckd���o���V�<z�u�*���o=of8�-�:�p���%����5p��(fC�}9��p�߼�mKd�6^� ���+��$������I#����+h��H��C��t�'�VI�,�J1 s;����r�8����sy��ק�����I���j�lG��h.`P}GM+�j9�g��a�C8�u���T�|N�e�,�vw=���2S����.h�بݛ6�<N�Q�<At�tq�)��5� S����C��u�Af�øC�����c��}m?�SU���Ƭ���ŭ�G"���.)�kp`5�>�����Rbm� 2$�#����ڞ��]Gsh�:�ň�Ano}�6�`JCW����`	�`���Ac'%�_�2߹����*�2�bN=z�;,@���i�'b��C��Z�?�aU��f���t����u3��.i|LlVQ�zc��"0�ܮڣ!��&?���7mQ����Vb�Tj4��)�=��P� �0vB�98�]:)�����"���y�hz���9m�P6{d�88��I������ k��x�h������6{�>�D)�� n=Pf������[K� 80���%�^⍭0@ć#�r���8�����_gj^v�<���ْy�mA&8����#����F���V�z*A��,(e�?_{Pb�T<��1��j�;���rUӲ�-ew�o�C�j��Wd9^�b	_D�岯l�9��²�l!4��jJ�f�l�+		k�V
�	���u=���b���ڟ�Q�y|#���H�]	f?�q�4I��P��z4i�%�)ސ��7���.����aS�LX�2;�����!<�љ��:[/:X7�1�⊄kM�K+,���o9pR�k��@�'�����S�y��߬�8��8xI[�����+ʥ�]�Dx�wӳ;��f+Dv?w0��Ö�����ȅ��ʄ��L��ǵ�峀��RL���s�`�i�]��AD�lg�ҩ��K�76��
"С����5�ֺ�[��|Il#:��»�����V��������i0�[en�\�&��?�x*��j~?�p��c���f�I�����7����00��/eJۻ��o_�O�d6?Ol6�af�w�����Q��-�ۃ{��5������`��H��3�x�i��^/���׶[RG�z�~2q���P�n�A�rh�����Gy]<��E���sJ$���<�N�"X��|����-�N�|�.�::G��J���M��g#�Ba*H��ޜ��_��8���^˼G+��m�~�ȿ�T����[�AM�� m��)m]_6����<�ɗJ�+��3}|������w��%C�FcFF �0�|?q���F-ف�1SA������R�R#�Y!��@oLb��K:h�޹���A���N2�E!l߅�d�k	ϟ�����2'��,5�S�;�vzj�҆�.�	o��t*�-�Ȑ��t�߭��ӊ��"?�}����A�mz�э%H����>�qj-��,���߄��`i��_#��,]�V��X������;��A`gS�S���-���`r�
Q��F4�e+�7�{���NX��G�@-���d�Ih�j�U:+�N
�f���[�e~��MZ���I�Y�������-���B�$���* ԁ-�~���솈���3�$�v*�<�4M,q͸o#�w� �B��,�t�)��Y�e!bO��9�E�(uᾘD'Lb������4�p�����A�`n��[��N���J �*�f���u�4�H��~:Xo�C�l)PC.���ס{�@�F�o������33J�+�O:B|V���f���o 7����i�����ޝ2DRj���ʛ"�>��7� p���N/R��o3�ݦ����pL1?XO�e-�p�֌��q_3��������bF� �;B�;�Z|�f�l����;�޶>'�Ed�	��S�G�����76w�}���5�+�Dm�yH�.d��F�h���K�Y�6�T��@��<a�5�W_@1����� r1Y?+��n���������������F�P���F�)����Pht��m��F�_ 5Or��.1{�%K�sҢ�ˏ�V���D/ ^����.Igy����J�DF�i��}Ls�fD��m^|�����FyzM�n3���e_=�k�j%!~!�t���>�����<�h���|V��n��MVF�(�/4wY��+��n�Ɨ��Sl�;�;��1�uQ��d\e`�~y����l]E5M����v������NfM����܃Z=��ˌ�x���e�g�,��b�IT�E���Yg�qH�W��z��\�>KZ�	ʽ뚰�*F��w������Nڼ�Pя��>Vk�����6����`s뚿x�<K
T�T�5k�)~C;���;���S>E�<}y���@
�ݭ��tӲ^;K
�Z��s�f�{3�TT���7]f��X�n���b���z�f�їP}��k$S��t���\���4Yl����j6)=2J&/&+�C?���v?�p3�~\D�zh ������bDD�?~���qa��sN�0��A[����r���RۙغگD���Ju7\,�2::�!�< �!A����y��T�.�x��"9�K�H��Y+��+F�L"FK����)�/y�/�K
?�������q$�"�"�EѸu��r��$�*x1t'ώs��H��>����[�iFͦ���W���Wl��`U��N5$5�'ڲ��'�����&��e�)U$�D2gM�=��x��4F�1̥]���?�{���ڶ~�$�ì2²��n�@�Q=�w���઀ycĵ�.�╄�[�<�f�.��8EЪoa��1����Wq.��Z�l�`Gg�N٪�TT���f��p"pv���i����ժ���6�4�oý�Y��1bVӬ�<�yq���v�1@Ê��wZz�:�VϏ��bL��j��y���Q�d����L�X��V	�`�#PU��p�o	������ۇ��L[�4��7K&D��ݿ���}�b�l��7NL��!�Uc�!2����C��^��6=`L�@5�"���8�������9�s�Jˉ���4��PoI�o�B�8�jџ�����l]u�g�{�^�q$�|���ޢ�Y���qP��F,�"��py�������o�%��4�Oz���g�e���c��t�IӴ{����1��H_�fͰ�L�	<i<hC�՗�f��H#��8�g�3�2��aEh~�D���!�9KyZeš��^���qWum�0�u4�j�5MA+��z������ף�m�8���#V������D3��9��+��7IG�k�X;W�&{�Ho���e׊�Cp����9�o���&wD�h�;��}���w�Μ��'P�ӕ�4�w��V�ؘ�|�**%�B� ��G�m���3�iy����,F�	�Y�;�@��F�$@E���� ���L3�\�LhlEa{Z
���e)�ꃟ EǏbau�H�!�	H�	��<��6�ج��4�Y���[�����{j��	�^]�=�s�Ov�l�4J��Ek��!X}?Td�yB�5����q�a6Ϋl���\�tY�<S9�J �_?�\�Us�V*R�����B��h�����p�si@C�SD�ns�@br�#����#R���z��"˚)��ݒkD�����K%���Yx8���6��gQh#o����?�#̺����^��ca�sVd�������sL��>$S�,O�n��f�3<f�S�2���/Or��ӌEk���`��P���\t˴G�$yx�q,�[��kAH<�d�v�}� B�W])��Ц�����ŉ�آ[����Z�C���\��|�)l�l�
HG3D�/����_�#��R��������������	�T�@u9����xaȜ	�Q�=�6�HO�	[AږT�R	�ai���e��I��%��g&��w�%�#��h_ǥ4�W�&�Bʖ��go {��%�y��aԜ������ ސ��L����	������i�b�v�I�k��M�qzC9�i,�#J�$�q�=�-�ө�������g,/���'�#f����"�6��F'�S2xw7H�k��O�/2�َ���E�k�x=�3x辅�?(��rޔr�=�25�9�١��%���mN�`6.2/q�Hev���7r��U�gDQ��4l4�z�q�����P��:㺚�4	B��U��?R��^�����P���{'W7��T�3���@k@_�L�o�|�~'�Ә�t�vd��Ļň�&��#���m�]��VC��C'#�J�g8�AsT^��TNe����m��rW�dP1B������゙�[���x��62Lae�h�����4�iRV�h{����Xkw|oh��i�M���LL��݈���'=�AXu�m����� G*Z���{��ER��*UW�u��̡+=����������^�-�w��}]<��ݿ'�Y]�y-¼g�[�u�s�lH]�#�	>�@r�=lb�r|�9�a�>Иi_��_�S�:,�E ךSd�0�d��<N�u�XU��p���d�/0yhr�R�aF���ISw�Bb�"㣗7���f��������,���u��E�X8(��.$a�n��Aږ��T9�����7?�q��Q�,�Jډ�Pk��+h�[ږCmI�����9��6�wF�2R<L<�K��^�{'�Foħ����A���w��-�Xs���\��VY��~���f�����<�U�]ϋv}�+�F8x���KYȋ>r����OwMs�5�t��R",F{s8��s��+	i8�)�m�i��;y�� '�d�:�֣�^]�
����V���z�0��ʘ��1�K��6�
vDi�.e��[�K��ϣ+�ي�R�Rq*4S�R��T�����O�k3OK��$XJdj�>��HW��8̀���"�k~q���@�4�O�X�t<�jB$q��g��v��/_���b�����|4��s&�|��k[�n��-�b
�u�A�k����I�|�jag#&�I8A"p�4�(�
ڋ�[�E&V0)�g��O�i讞��<k�)A/�z���'��j��h�s`��('K���!GYS<QA��b	�}��	�칡/�¶5G�?@d���q����~���ԥ�3��p}���_�Ò�e��޵�l�M4�1�f}U�cA������th3(��0I;upbϲ���\����4#�!#��)���7���I����}��x�V*�2����T(Z_v�q����O�d|�9_v����̿�f�n�+D*(1���)Q{�ao���%�W*���H�Ð{<��v�,�n$�V��;p{�6 SB{�|<f�Y0YTXB��ܪ� 꾵���4[KD4�Nc?#Cx0�W�ZZU�O�x��E�6�)�4b���b
͖V�w�=��Q�5ٸ�0�"�O�@�Ak�i����z[զ;:t	��@��S|g�I���j���� �㓅�>lcR,�e4j��<!��|D_|�Z�%��2�C��dL��Z鍽!�d�V�)Y�A޹gƚ�%� 4�
��5@5䨺�����&�=�C�[���0�0j��x>�+�:��k� �mLB�lD�K�2uu� [09|򨰛EƸB�P�����O��$\f	S�s��\��x�`����So-yj��`q��ڻ(��V@Q�R���0SJTdZkX�y��%����=m�����"��W0�HN@�Q0c�����rN*MMCB+���#�m�<R���D�R��%լ���M��n�EՈ�vI�޹�D�H��Y V�/��[٧��-O-��[��K-��/p��%�7�hĬ��"�j5�����:�R����O�o/�/f��A���qP���E!2a*C�0��I�����XwG8�5��e3/��@�Z��.$]^b������2B�<��	&#�0[�����Ϸ	򆨦\�ݡ�Y�6 BX-s��ٳ�U�cvN� �'��!���R;|eqZ7���m���x-U�5%#��.r��_�i��lY���.��$m0>��)e��	�Q�q?`E0�3��0*�ܓ�Fb�t�#!-�'�Ǩ)���$��`���	�$p9�i.%VOY"X[�;t�`̗��:�X�)E�,�Y:e'��+)�Ȗ�'o�1Dٲ^���[� �֧�76�����ă���1������}�����J}�[�m]k��X����u��ߢL����H��)�� VR�D�Ш�`�\�N��#�I�j��=�m����L7����T$��}��!u[��(Bk%�����Apŗ��n�D������6(b�f�"�M$p�.�!�(�P|~$j0QNBV���e���隐F�wZ��{u������}�[y�=X+���CQX�Î9
0ɍ�&UZu]Iג6��+��GS��34�I2 z�)��2j3�^N��
 ծOğ�HIRV����ؘ���l0�/c٦�:N_仅3���-�z���畽������(��*j2�[L�ab3X�Ѥ�z�F3_Z�����:'�%��ϼ�S�[�������8�ɼ��?��:�m��M�Q���V��n�d�ؠhr��#��U��
(5�>�y�g¦	V�@�.E���Q!��F}�F�|.�\I˾���O%*�?��E}v��9�N���I���#���E��7ڞʓ��9����V�W��{*�zj�\�a�-�B�1�uV�8�G'mH���W�ˡ�5�R>�N��|�Db'��bQ�]��`nP�0)�b#:Ok{�B�6Y|eɰ�ռ�O@��KK#�b F2�e`��پ�JK�Ͱa�-���ȭ_�h�*�N�����E�a'�U�;���ǆЫbE��d���;�8���\j��7�QN����%��:��f��K�� �2������Z���`'<61�&=�}�G�c3���L�!���4�@|�H�5��9?�4��D������u���4��|C���&���q�ԅ��l���pZ���W�����EQ틜C�;�7j��/�EI:���o����F�(T;1���H+Q�]~�k�ǐ<F-ݬ�S�hK�{Y�p��Vo�%7�]A�p�����x��4)�!ϱ�d��?/N�%j, <Ѵ���r���g��y��N��?S���la���J��`f�-XF�:~�Cg�~��nO[�4��U���� ��/r(�uLKư��a��P�JT�cp�j�A/��C���j�0!���|�"!���"&>B�� ��o)
����jC��"�í�ri�8���-R'\�5���k�i�p{��𣱺�����)V���H��1f7p����Wf�E�c��6��+X�9ŒE$�͞�
�N-釣��p�fp�?�T�AS�J�m�]#����P�� Utl }��7c*��u^h�U�U@haMc\D�f�-`"�L��+�א�B+����50� �_!�C��,U�O�ysWI�$�7�6��rտ�~?V����n��������l�������"�[�\v3���H�&�}��bN&_F}��x`="쉼����o+��\�ʨ~T��Z�)g9��ʆ�@��$	��`��r�}��/��[\t�!���~�~\V7��Q�h��%��E�݅/�0��v;��,Nߜ�V�P��LG~-~������R�y�P>�ۯ���5�C�s����$M�ٜB��N�E ��!t����� ���-�t�רh��5�|AU߂�θ=�	"�ų >�^����(?�]����Bg�f�lhGR���aN��}+	U���������/lD�I��Y�P*,��H�h�i�T���|�A$��ܙ߷�i�B^/����#�|Z����C�	�%}Չ,cbeKBy ����T����bf{�o��Vѿ�q2&+�s�av��r������ 5s[O�A7���lI�:2e�`!�2ڏ�A�	x}���GY��ka���ǎW;ۺ�[�Zg�z�PR��L�*vS�gx2n��b,�n�08��'��ځϽ7���K�3�!�-��jn���Hip��iځ�. ���R��b{�VB������3�3u%��c���}���')S�d�¾Q����mYt���걐̏����LN,I�t�76����'$�<@��J�y)��h��Z��A�F������/��~�#��I�Of���]�A�#\@<߉�pm�V�?��X7�����'�L���� F �+�k�9�6�q~W����#櫷&%z�:V�5�0�KF�̡X?�R9�3�9asY_Ǽ_O��~�iҪa�i`v�%�#T:�����9��m��8Q�k?��Y�#E��2c��f���znR��]W�V~c�J�i�i�O���F������LG��r�O�{a^�$I� ��<�(����F�����}�h�F��q��HM��A�/L����$���^V��G):i�]���+��*�}���a=ϛ�Ő�UKɞm�	P��(�ج�0}�#s�H�]%髒f�i�����r��&-�@���U������\gD̘z����G�����<��#O��q��W��=0��|�h*��>��(���+�l�:G�59!�𘣎 a*��n,&~�T����_ ��1 ax1�(W֓�>���Ih��	�Z���A����zD�B���黳��͂@�	�k#��9�!� ]����$�?��E��3F�o<YV��6�W�M:q��,�B��'\�0�j�����XH��(�������/���16�V��H��(R:sk��i�
�(u��Z��8Ӧ�/`�VUT+�@-���H�UYr�Q�?�rW9k[7
�A�n��j�>�4�~� ~b�>t����@���[[� �,�@#�(��`E�g2h�m��W��d�7p�J\bCTUZ����jQ�4L��f���g��	����q� �!�#�9���e����8"^��R���[M���!���A]�=����j���T��l�N�2���IK1�UV� �d�|P�g��bه�?�m��/�������[�:t�/�Y��|bV�?b0Ϯu޸V�L������mo�}���,�1���������TCHA��5tW�&�D�e�y{+��M�T s��)
�o����@�
b6a�4'Tܬ=�Vk�J��Q0�~^zcR-Ѽ�(+M�JPO�J7�X0w\qT�Mnj��Z�$�y�D؋����'Eh�@��r����tv�0�h�(������ɣ�J`�z�����}%x��HX�[,��`�ߧ�-#m���Dd���h�Fe��"���rY���X��% �u���(�$�J��y��v*�o@ +����\(�1������	
�ֻ$�����4y}��*i��	�r'F�Q��]�o.�92��$��r��y[�C>%�@$4�L>"��E(�|�]��$�\5 ~����vDs��O�7c6m�vŎ#�9�w�{ �������`�w�;aK|��u���%�������?S�Ni�ңЏo�QS�=��hbq�K% � K�֍S��r�Ø��I�mCLKz:�Gr2�o��y���z��#�_�`����{�ِ#/�8'X�m����O0*�h��ܜu�t�b#'P�7��0�#�@d���v����pif6��Z���k!V4(�°��p����O���R�甐{
_aE�@��<-�X��M�C�*fy	7]O87t�h���;ĈR��>�,�Q?ٽT46JXx��)O�4�
�'�=
jv�k6ͱ.��˓�����B 3sVM�_��geh���Z��!#f�08�᜝#r=�45��Bm��8��Ic���v̰sd�i��&O⧻3�^���_���J�n�н������n�a�eS� ��^��+O�J��s �ɟfzx��%7����
_-�&�$�u�^p<�R)����^K�}6�*��`Rꥥ㫹u|"�f�=%i�A�Pp���Y�9�I{rB̢5!����f��z�"O}�"UXvi����prMb��X���5���i��s��ሤP�`��t9�x'���Sq�Wg�:E�6`�p�Z+[ώ*B"?=M��rs���!�8z�Ȉ�5�]��J�a/Gr�3��ASq�f�V�e�o��EƩ��(N�-r�(Km��m���8�������N���O��<����^Fv�a�`V�5�<�ɽ. 2�SOx�G �WhD�����L�(���L"p�i�O�q�^��~B\��΀��KH���O�F'=�\�y��2�~�J{�!�f����;l:b�Oڦo��ԑ�����>Z�d��{����$��똺�$�8<MD}��\�,S�P�$n�>ɣ����K�+gb�� Ojݐq*E��W��"0W,%fc�n��Le�J�f���(����3�3�p����!2�拮`=�������i�D8BLMy�wę
'�V�Y�����iHE��x�����	0�ʒ�L���ǜU��G)*V�i��f�D�!��8ѕ� �d�9�Ybv-x/��}����c��S69�~"60-���YkC���Ǌ�Y4�Ns�N�A�J꩜���q�έ�q�_���<P��e|S��)z^&�z	��v�gR�����T�.p�� �/�y�D3�E�BY=�{e�ZD�9ǩ�v�|1��]���2.�m�3�FE��Z\&T��BoY�����n6����o�3vv�j���K3�A�\S޺}��? ĥ=p�䖋��ԯ����o�5 /����H#m��"���=��k+�S� o�-�bʢ��K�`<��2#H�k'�8��A��pH��_k�D}��	!�U��qL\E�~�nA§�̵�&F(D�2��uO�h��~�C;=�C�M�ݱ���h�T�Fųł�^n����7�A���bd��]E�ք�ʓ��!+�$]ʸ��w4ˈ0�B�Ub�ҚW���W�3�٩���B����Z+�#,�Q�S#��$<jjI�Ko�k����搙tH�Q���v��:3�/��Z��� �m�P/}��v��rCz��TcV[�T��G�עU�*NL���'�Q�K��/-��#�� ��\��ݽg�����|�o�l0�Zb__�x�.w��؉h��������f�b��qi �Q�ݼ�Y%�D`<�O��h���jS��%�X��C~r��5o�X�.���H�c'�v��ڮ8�" '��� �B����5��t`*�N�8V�s�����D�]�)A��@�>�
�^���ec����\#�έ�����j��CW�{����$/ȹt��s� ���%E�_�|�W�0�/������p�̇�B}�`<w�����e�k��7hKF���$yA���|��ᖭ��NYq�4�"\���	G�Xtmy^g��/�Ё1�M.˱>C��S/7��;��ri�?N�{[J�� �GU�$�)���Vq��;(j��5�ᮣ6gqOf��D�N�[a홫zQ1���Ĕ����R	�~>D3�������L`�F^��;��vz{ǳ}��Ɏ�j/��W���}�o����xr����+��]v>�w�W *!��b!Y{BU̽
]���h@����%ɕ$�C��}&q�W��s0z�r�h��@�v_�f1��ƴ*(m�Ϻ5��F�)i�m@d� �����ެ��d�`�o���(��.�A@�V\�ƭx���f(�c�cp���	�P~�d�1��*����Z	Ҩ�/�ﳃ�0~ySI
��Cc
����#`8un�����~�Û�4��a�8>���u��dT��s��T�rf�bMV�F�\n���!�`��N�k��+Sֿ���|�Y���k�xYo��8�;)�N�� ��SVT#�)]qD�!�U�HH�B�8o�������fG�����肖�-ް����[6�P0�֤�Zr����+3Y������C�����'�_.�7N��,!��Jg�1��+�ca�l<�5��kĞ�d���W�]�V0S���Bw�'��Չ�,�x[�\`VG	^$L�*a?v'il�W�F?�Uqbi�z 9���u���/�����;^�I�&�'���=��>�<`!�V}p����=�G���fd��3��]G7$�i���.�B8�Q�Ɓ2Ŵ�ȸ;�g��h��Ї'��bў�,B��\��`덫x,&7RQ�h��ۣ�=�u��z�J��$zi���	/2��4�9&j��_�ȁ�->X,�u����6C�Z�n.�v����w��e?��:��`�<`3ޣ��R�9dJfc�cu����q���	��~j��2�.�c�v��qe��,Ą�B� Q������C��jw߶@׮f2���?{�+d��yq��i�B���I��K�b*�aHX>�8��!8�:�4ў����T⾸F�y�veܨ�4�i綱�c�����d�$�b�������yvr�ӄ�J�缁�3,J�q�k�����zX������f�#�Օ';s!+���_�q���r�'���*��9��qT��x�@a1a�v�^�@�jGSూ�J��k ��I�ت���������IO�*g�|sߠ� p�Q�����Lj���T��1���[MD\��If���~1�[�t�Q<7����5��h��8�h
K1�6��Hn��Jh�3�x��m��&U��� x��� ô��8�i5��w�o1}����~�sݯ_a�:��iG�\
�;CJӌ��t��Gl:_��O��R���2?����������4��Yπz�s7·	� i����[{c����t�JU>�vn�+�v6��K�6*��}��O򺡺�)d!NV�NՉ���Yk��I��S���LX���jk:'Y��أ KW�x�i���nKI�
 �2)��=�����N}&�\Onʶ�a!Ќ�!6�-�{H���Z`x `�e�as���jąH'��b���X�k���]�jP��w�M-L����� -�z�m`ƣZ&�~k�?,�$���������ɧ��+�����=��@�� _�m���TըK�2"ὦ��Z�=KJBq�~��z�E�;0w���k56��i}���1�BA���c�R�����`t��ڕ�>WkY.\I�ڪ��2T�w�[�� �<!�z���W�_�u�:�S�|x�7�"K��C���SAn�o��wЬsMK�����Hm��1�ǂ�ՐC�>n!�;,T�\2�E�],k%�H\����4-��������5�?8���a?�A�)@F8wtt����M|.�A,p/��ڜ�|��:О�Ǭ�QRuu�V��<V)��]��w�ްĨ�CR}1t)��9���s��?:��/� �Sj:	햼�s��.ܛ���ߑ��p�[��:��)s,�V�R�����o������&��z0.A�U[l�%���@l�䠣\;���ɗ3}�8�t���r�=�k�s�o&�
���o�0y1aP����ƽ7��S)dΦ���25 ՑM��vg�����D��uSh���>)�9�ui~�x��VR���''uc��n	�6��߽��La#O�s�(�(���<��&��Uϛ̸G�U�m&�>����gl��͝{�[�cx�7����|c��Gn�5���9�w��-�]���3S�=�g}k�C!=�ī�!z���X����r�ύ�Iۊ�Y4�Fjt܉�W��>�C!-'��
e�0�������/�eg֙�e z!xSm�7E��f}��[ﴑ]�3\@�_��C������î������ffmuמB~���ҹ�E���OV�kWJ%0Z_��
� O|P`E1�6��y���RP��}U�����d�ðWn£�eIf��&�,��{��"�z�5I�e��*m��y7�MNkT��^�ֈ	J����ry����ǃ7$�O�k��+�k5#'�\~WՌm�9S"b���$��J�~f��,D��I�%�P N6��e*è�J~!_ɭ�%�h�
>̄����m����j���U[�}�gg�( /�_q��k:Nw�jq�t���`J�xY���@,�l����F�+�[�0�5bx A�fv����8����K�٧W��^�����\.��c�o��k�R��-�7���%Q�cR4<YVm	��O�E(��I�z�5��@|���u��|�%�鋫8^�
d�$���f7ʈ=x�"�kPd�r�k=�A֗�j
"a�  {��%)}��A��1�����%s$��I��� ���?�с5�m�&�~(y,�z~7N9�+2�㻈��	b]S�3E\MQ����*B��z�{�{c9�����69y�t�]�N�k�-��U^���R����M��;2�T݀A>c'�e���S���)�����y�p�V,�� �G�KC�b&W^D�P�
�8ب��E�`��^����|�G�Ӛ,�p�鞙��ocHƍ��
��=���`m�0�
O��.2���&9�o���3P4�d*VEM�]�������e�\�d (��jQ�����<O$�)\` �����|�����@8��c AHov�X��3K_�����ʶ�����K��Y�������������Nt����*T� ��7�x��Vu2I�h~����zTR�[��O475�??d�p�~����u%ڰ{s1(�?�����I>���Y(P�L7��NG`�X��Cʣ;<Q`+�$d��Q=���5<d4^���M(�b}a\B�h'^2���ڻ��v��򅻻7�ջ�� ��rţ��X����1ՐÛ���b\ڛ3k7k~q��FP<�ퟷX�'�ߘ� yD9rVQp��(I���&��@�L;L�V=�r��5�d��2�Y�H����*Ex�3����QzaBcj�r�w{�k1��{�_4y���"����q�����V�S-�%Ǔ�H� S���?�~��ן �۸���Ţ�) �e�Lr~a���2c�_�o�Oe])�����t��Ϊȼ�,1E�~ �WvȐ�*G�iyп�%D�g�';䭞�B��N�G���_���N<�����G��yt���r�W�ku;\6�@���.��戩�����i}$�x��Xp$�]�y�r&0}�Y}>���h�)9�e���A�6���sw���eA}9��wu��8��H�^�3�Bwad�d�% U#�Bmo��j��;�W+���
׾�f�w������!�3���C$F^^���(���#f�]������i���S��������No���_1�B���i3w��u�aH��I�G�,w�R1��&8wKc�Bp��;SA|:�T.D��d@�@���
��?�A�&��Z�?�,��Mn��>�� ��z��O.ƛg���y�`�0K�{;Ht��84lV�V��n��?�?0�T��ھ�J�W2ca�sa��|���t�n�iOj�V��Na�̰�������K�B�
�܁��7]����Y*��+=��ۙ�b��9�9���������$��B�fa�Ū��nO�����=ȭ��'��v=~G	���Jˏ��C��L��.��=�2R���������� �$����M�d!��cw1�{}q0�wxV��i��C�t"Ł)����G��U����#��.�����+��LS^V�j�r�'L鯲���D�M3D["b����@K�T�ak��/$ܽ��A^ X����t�G�2`s���<��7:��w�NζFF����r��I�>�H�n��vS����˴(�T��95:&�a[U�Z� 3�}L��5���@^��"x����%f�M����}�c�#d7�0�|�
�)i���S�b�-�v��[C�yS uEDޔ�6�Q�ż����+���q�$/@Q@|�Tt:r7`��>=��3$��".�#���J�dk��N`<����Y'��a�+�Qdo�,�i�B�8%��`y���Ju"�v����^�]!?
"Հ���S����åG�0z2�N�{Xm��
�'�~v`D�6p��IP�F��j�����eǈ$�l~"#�>0����CS�oF�����v�Ư�!��.𙬥�wV� _�D�G;�t�����.�QF7�XWLG	�8�y�?��Z�_n����:j��F��i�2�p�S�h٬�K�7���q�I]cƍ��B�tf������']�웅�C����S|�U�gy1gwI��
l���ĉ��[X�-�+�w�R�I4q/���U���E���T���!0Q�U�=шү�)�<:�<x��[��*s��໌�#��شc�E��X����M��.��eR^��8�Z���k3aR��u铙�V���'{���k(
f�����e�;��;��I��:�^O�1�c0�
M�)J���n�8[����x�O��e��k4tK��⮶���ڂ|tW�0zfđS��A������$cjW�y�6�@��h$��{�}QM{c|A�࡬3��lqeoZs�Gj���a�=�t��'��"��;�њ�D�q{��ț᱗a�,M���PEA7���ρ�aO	�����	�ۤ�*k�b�w���t�M��6�鵪O*)<�F�҄+O��~�uE�OX��A�j�ʪ&�+��&�J�zP��H�怳V������<Zd�"�ז���	f��"��6Eoa��H�!7�&�Ǯ}]��������&�;Q>�������d4�)�u�`�7=T����/�=Ų����[���ng�g���k�p�X���G�/��i2E�^����Lk�v*�Z91̦1;����6'�/*������K+��SM��NL� �e��$����BR7u��j'gJ���S`��R�\�,bE�L���B���ޟ�55�	�?�Zx�^}���ʭZ&�p������Hi�ּ� ����^��sC+���A�h>�;�5�ʷ��u�w�!��A)�m��(�	1�Ugkˍh��!Z #�U��2�R��fWMFwU�n�8[��'-8��t�Ƚ|�jI�<ǭ`��?	&�	/[5�b��Ѳ-�kc/lmDU>�cp�"@����y=^	@uy��I��UڙM��n�bM�3�F�ێ�Z��K�.*���a��޾�YIxn�c��<o���˶�v	�u��*�E��A�ZWI�~Ho`��y�m����%�#��ef�����FE%�b���A��i�a�������������8նqv�~�`e\_���>��|e�5ꢫ���ޅ���h������>�(� û�# #�ʲ|�)`�y����j2ƛl
�)3�x��;��h��
	I{G�1�QǳhX(�Nί��9�C�#�R9�Np�!�XHs)�Ϫ��� z'��ήI�[���t�('>̆j����I;�`B�K>[\��J7�ZO��\��.�,���)p�KʈyO���@@��o�v�_�\�<t�ҋ3������+���n�D�S�e!䛦��E�����ك;f���,����i��o�헉�1|�Nƨ��6Ż�3���zi��h��Z��m-x�f2%i����pV�&��5����੷3P.��`%��7�0��y�8K�F5�?�<	֏���
�/����ϣ�1�c곾7�'&�[&)�C�\%���R�t�`��"$��#�x��C�����̯��e��o�q��R�
�7?��5�7L������LOX_exub�Sg��EZ]D����%�-�%�����Oۋ�s���Ӧ�����ep�7c�J#Ҽ0��4x�3g�P툄��p/�o+��C��O��m���i�3bn�5T��G��{��i �(������sS���ʹ���@Th;�&n ��|5x{�#ӂ�E�@�~H-�=8g7�tA���}![n/{-Y�Ō�r:Yp�Z�U��0��ǿ2��\Av�.X%�et����o93��$T�#K�e�4q��ti�k�-��)�lgH��:�ǀ�2��[[6ۦ���md���\��*5�>��hT�Ǭ�ء���@�3Sq��$���e�ž._���^��@��e��u%Loh� }����Ss�\,1F�1�>�!'QM�I�c�ꮥey<��F��������r PfaJ�d�>���T�#��k_����4l��!#Lk�Ͱ��S�<����=92�P����_�5�E�����[A:�G��(�KB9�&���;@.�`t\jo���o:a����?I�z$��l��4�g��{;a����6�¨�x��0��.8{{��x��A��Nڥ�����S�q�F�BT.��"&�"L���ƫ@	�ٽ�(T�B�>�+򑋳��?-HYs���"����R)�>��v<ѕZ@����T59Z�Ǉ2X�"�u��r�@��s�];;@�H��������r���}x,�GK)��臙e}�CuZ�F�K�s�J=�f! �8��e�朩�/bU�Jَ8�P�L��f�gkB�9#z�$F%��5w6ȪA+�4q�c'��v79��4��p�e ���B��l�m��BV8���`�˛�	�oG�����uqR����:t���Я ��p���U�N�̇U�je�!K�|�4h4R�i�)��ɓp���(q�k���#{��VŃ�X��^��=�s*_�>��ƪ��1,�{��EA)�Vn�c����ȱ|�!�&h]�h,3�v�6���	OC���ډLs�DJ��T���K�	/�<���P�K(�ߺ��ܖ������^>C�����_^E��i������9��7�}��i�[7$�M��a�s���#��60T�'�aAH@d��8���@�	n����W��"�*[<��E`����&�R���7���-+��gFa�A�K���B[v�l4�кA�-�d&\���S蓹��$3)�y������}	�)v���4"���4I�� ����U���L�?�q=���}��(=UC�"r�!^�1�SMH�q�x	�4�͛�&�wn�sC��G��芣]M1O��L�����ĕ������OH�$ā����j�z�H���}�A�������*�LRR�k��߂6���6����UU����Ⱦ��A��Q4K�4a+��᧼�'��@T8�.��7�{��q4:�sd@g�g�>�Q����K��`�� �/����Z��M>��&x�&��w4���;s����>��y�,��&�g�ֻ0Ń�9���n�����0[�fL��M�(�����C��<����Ę^>COs�ğ�n[e�yx�|� ��V�NC��)�����ꯊ����B4��"�h�K\����+)��0�P8�xF��0�K��")R�'�&]�3�����+y��ͅ^�,�n���p��ۣ�����y��U�����T���]�_�)9��y��`��W�E�Z�1�����%4x��HM����Qғ���P���;�q��6�<��s������;&/z�!-9ݑ��:Ip��c�D�4�Y��G�Ei ��f(�� e��Ak�VQvl'�;����M��?�m�\[)rIc�\C�ů�2��x��
��G�!cF��?3J���oN�_��!��������6�v��Ac�,�h��Y���q$>�O 1	��z�7پ���T�2���E1Z���M;��?���W�gC��r'���p�_)��>��b��7 ��cj�J�wjY�[���}��5n^�e2$tZw4�A�b\������g��L�4ŲD0��@�<.�<�9ރ4phOCC��Xbv��f�V������ə8��[�^�Q��k���=ys�l�RSL��>�s0�KL�|pd54c����
�"��so1��2�oo+����w�[������y8�`�� ���|��Z�l��"�b�V�_wFu�<퀔�5�2��{���W�A�`Gр/c}P����y���R���+ܟ�k�Ib�)���b�&�����Q/�7�9�j|f��fA�R,��s5*��'�E Z�N�K��Q���E}}�f��e�@��,�����$�r.���siK�̮HI�'	7iq-'�}��,Ԭ��̢���&��1!O���t�S��q���\�+��yʯ�"��q'��bO���}R*ک�N�v�u��p{�y���糄k��p՗m�àJg���rz���d{7W�ĚO-+��a���BVR�I�Y��s�h��)��u
��gs��gMc�9�z���CSI��
Q�J�z�~����D-b��k%[���*�t��|N����f�uJwwd����s�M<���o;r~{E#����{��~9��=���B�7�4��	G�~}�ؖm]����]ݴ�nn��F~I*���tE�5��,���(���6�S�
=u���Ja�0�=OV?ҀH�?be6BR�d���D��U�J�� ��\�^�4m)�x[!57���~����fwv��+��]���D^��;Z�dP�Jq�_J���gf���=���]���n۽���{��Al~&؇q���Fy�~!���>͝�;��2�e�n[|ت����Wf�L6�b<�:�%��|��*�צ�������-ve3q�M�.�k��O`�9�� Z윦�2}^iD64[�@��w:G� /FrZ*V��(���s�f�֘�֞
Q���1�����{�Z�W�sHLf�!���H�����*���M	5h�|=��G�O����7Y[�r��&�י+rE��v������T��$��,xó��n���-	��vOo7 >�a�����%P_�0�+Mc+�Ƥ�.NaW]G]u�p�d�x�n���GS��" 71e�1J�`o�C�"y
2��P�Ό��G	ܦ
=S�G�%�>��{������5�U�޽T0vn�y{�}����AB�d��+�w˛n�~ܼ�{������x_�A߳K֪���\'��a\|��T7�kW�y�^.��:+3ڂ,�o���k��Á��9V5�	Q杁A�M�g�x�9X#	��,�����Bg���cL�[�y�|qD��� 8�(+�7c-���MW[���(?�V��6�I�^�`����w�	���-��N�m'T^#0��T��[ݶ�����~�8�r�t�;� 1B��|w�^9��3��s�	֯��|�<���Y��!\�C��R���I���;�}I�━�VHF�YQ�L$�H����	�L��xK^b�`�Ŀ=�C<�,����.W��JFa`,7�g,	��h��� $zSsj�`;P�#~�h����c�"����S��Rl����b�:��-�M͸L˪�L�Y;p��B���<aw~�r7���\�N�;V'����C����قY >0���P4��N9� �g��\j3��s:�I��-.�������_����۳`x�A����
�{��ޤ�׾���j�OMƯ�:ݎ�<�r����3��q`�[�\��"��5�E�n��F��@��"�d�_���mA9}�'*j��U��k�s�6��d��� w��F��Vtp�!Vy5N����1I������� ����G��_�ވF4V�x�$9̰`�1d��@0��f��^��l,D��}��(�}�,��<=S`v�4�c��ru���S�W���u|L��6��CbYɈ[l��ҥ��ޭՒ0���:.�-7�<�D�K^J=0L�� p(��\�Q�&$���B[l�d��%�Cj/Ȁ��Y*�j�Tَ�ȟ��˟��8\֯��ۆ�d�tAf�+�<�����
=��{�O���r���#��(�3	'!R~�&���
? �Sa?�Ms��J,��iD5�j�u���Z�Qu"6��%��[��X��~�Td� ���u�,E�+�21f($�����s�U���ҍ�r}�=fpq�v��>A�v�hE"�5Ƚi�y����x&�gj�|�%1��}F�EF��U��E}z�"��|����(E=
�+�?8�����_�#*�tQ֍���ѝG�Ub^��\��Ϥ^�3zE�=Q�z��9L��B�V״��c�)9<��Ǭ4��L�Ks��Ͼ򬇶'xn��WZ�1������q7���!���L<��@>��I^�)ۜ�[�d�\l����-]#��?�����g�e�_�zig�9�F���Tt�6�t����{sGca�5$O ^aa)�l�������΁����8�Ӗ��@_-v��u�6<;�钗al�'�ص&:�q,Y�tKVg�ĳc��qm�Hs/��/�?5:���Qed,�s��rTuG:)s]vh�	�-�т��B�(������j��4�-�玲q����:�<w������	k��?Y�
`x�����x��c*����O!�E+nաx�mW�dh�=e�hҨ��H�Uq+��
�b���N�����O|̵�J>�αJd��Xeb�z�%�Rc�<���$����k�Ko�QD?�od(@5 ��0G>01u&�%i�Fc��*ʸ3k�ؤ_�~���~�^��(�ζ�O�~(�K[��~+�Ћ�U�g9��UD�����d�dB�^���a��Zc�ۦB\�a��ޒ��{�%��R������}_֡c��O��c�[�8�xP�c|gxrR��`��B���p1`P���I�os���4�~��"BW<g�a[��OQ�g�ݒ1Tz���S?|[�X�a�8����y�0t�5Ձ(H7D,j{]j����3j$,����kD�[U�'XdZV���_8N3�e�^/�h��X�HJ�ːa��ڽK�^T�Fi*�)�-ҿFw�7��9Cn���GX\�G
!p��cx��P5؟����ZX^z_}X7�h\��[8�����:��i&��o�/��~��د�,��8�[ס,ښ�TĨϒO���y���gl�A��!L��U-Zc�%�"�sif[X���q i�����~�g�U� ��rF���:��H�T���!x/�F��x��0�K�Q#f�ok�*������m��0�p�*3s{�^��,|�K�I��5Wʊ��U.�ch��t�+��	���|(N����&���T���>g�n�(3ѣ�G���9�����7���[J#��>|j!�\����Dx�;���Sn�����KD��6	]���h�:�W�v�S�,�Ϝ��Ҿ�tT)V����+JS�!�`w}7��=�z��¬3�˳/Rǒ�K�,�,pO�<���wRp�˹ͥ
��!�g6�a�rC>Hl_�����!b�
^�`!�J}Y7�%	p�a���E��	o%�S�6T**C��98�;�8�j�����<b�ގ��T$����0��>g��n�=M�/�$&��T��<��6-jN���H'���X����z����:����>h���o�@�����k,��Q"��&����?��0v���yd`]�SHMq�+���r��Yg���q��P��LH��Z�5����������dJ��3�'wS�Kp�g;���h�-�U�!�����q����4�����'8ؽo ����??	]�u'�*->������+Q"�JIV���hW\�e@-{�G�������3c'��T
�bl2m&���V��qp�L%\��?e����t���9�is�_ͪݮ㑝<Vcha7>%U��
q���TN־ ��7�ʶ��!g�"a^�2Y�7��S�H��!&U�G������ڝ�A�^�S�UV���e�-T\#s���8�Y0����=������[�$��� �/{RE����.����4~I�_����I��;�d����Ԑ�-�0԰5 h(�Տ&�����D�'*Sʻ�t��a�,�,����3���i=;��G�_u염"�c;5E���-��Kǩ�иj�#�4	�"�����P+�k:�h��arN���P��q"�X��><o���T��҅	�n��ɒxV�QHV/��$�eN5�~�#d�Y��M���P;�v�>y�GO�����S$t$��d$��jdc�gnD~[�B�7�n�M�gHq6or��q��4�#��r�bE�Į~�e9ƞ-�w�QUw|��$�zVJ[���;2J���?�� �;R�O�������O�`dIE��� �2jY_H)�{���A��lM��5��p*��I^;9�}�.�2sa��98�+�V
��9�E��e��*��-fY{R��Q���N$&�w���86T����u�|҅�ì�>#�__:�:���,��^��o�`h���qC(1(`���	��<��g�P�������\9��*Dz�)�A�<�u��6�v/�=XIKLS��C3��,h�S�+ �A"R$ˮ��ۣ����h��yWI�Ւh�B(��f��FbJ����0J!-^f���ԆA�"�K*�@�E^�24"�����17���gKP����$(L!�Y�j�H�ŇA�ߣB�*�$&|
@1��fGC�SQ��*lڙ�R~��=6\�X�/Q��y��[�Mݳ�#l	���u���+@�� �'��g/�8�Z�i��#�<k�Ze��d��P���7{-�|��lJ-Z���<`�\g4|�b�����Y�9�:kң�zN.�T+
[d�[|�.�I1(y���)U������oY�1�}��ty!@��t�N����S�y�ʦ-�ū�W�����M./[L�Y�;��8�$r݋y�x8D���{�7�á���+e��Ѹ���G̐i���6����^��i�6
�D7��3��	;w�N�\Ȫһ�Nx7
����	s�S�a=�͛v�}�(�b�����-���'8*nv&|�:sd����g�w���
ҧeԶP���2O��Sh�O���
���j�V��'�������Y�P�o���4ۭ�Ѣ�+[�_	`@��܇0��\��!�ו簪�ϵ�y1UŬQ��Tov�>xҒIz����c~�b� _&/�d�j8���/73�7�P���%4��EϦ�P�O��%��.?�?7-\/�x��k0��L�XU��rX�f<�~T�׎��Aq,�����pM�̀wԁg]f�Xُ#�徆��5�A_;��jG�׫3�t
 �{S�<t�S��"%ѩ���!ʵ�j<����n5���E2��7�q�{F��I�����UF9���ߌ_A�
:��V&�#��		�K%�X�4�_@�7 ��_9ȫH�)_���lvX�_�L��H��믏�q`��M�o�/.��R����9�G�U8/i��6���t��ܱ��z�'�C[�������ZF�I�}cM�mŬ��V ���Z��8���[1���YV��#������*�a ��Ƅ�]�q.����A����0�Z��ꋦ`Р�������s�{:�l���d��'Ǯ �I��W3��n�i�:�Ԋ�&�Hi��~��Z,��]���bh���_���Ju(2���z����t����{�"WyU46����]�H����Ak{ %7������}�b��&fV���]��xE0�;�s,o���y�'��Vu�ڱ��˭S�o���:I�k�o�7G0��'��'��V�{�V�^r�`�����$���
��&�&�Y�du�@,F��l\���AZc��<R���$�����]�A<4%�zاT����ӏ��C��w^����p)�v!{~
F��n؅�q�.r&&[�Ez��.L$��������pSB��ߚ:;�X�bz�,Ƀ�{t�@�Ee�V7� �ֻ6�C �MN]��*�L̜�����dE�}��`#罿�m��K:�l� �k͡üTD�!}l�N���ɗ���y�b��w>YF�5	] ط-����+-�⬟S2;�n$���~)]�V�ꔕ�o�'pC$���N�)6�{N�~AZZů٤ֻ�W��&}|D��`��wEЌ���n��]*szt��b�A����\S��YHuD����EU��I����o���'��	��$�+��ԼF���vYM!f�j:����!�Ãu�M��>��OR��%�x��oW�������,��\���׾〣8�.��QƩ'Ըx���7�I��."�y%�
�G_��
���P*�����@���C_4�
ӽqz����X���s���^��y��2����PR�ݯRWW����j[D��M�Sᵩ��,a�|�T�JٛwK�фӤ�)����m�
${Զ�{����`�,���B�= ��<�5��xa im �>�#�Cd�`�.��G����U�Ս9��N5�Bl>yf��2 ��������-�� �U�G��E���w��4_���iܙL�bfc��=�{����ә��O�З�C>_R/Q�0��2�N��*�C	F��
R=�ZB��_�FlU��4!z�+[���G�#���Vqk] �ئ�l�=;/���%j���_o�7����5?�\���k �� ��[s����i�`"Oz��|Ɯ�]$W��0��&����4�޿��WҠ5�Ŝ]�)2KY�E7t�%�mO�1l�����ǀz�V�@\�w�c[QU�Z���`�?�";��K�8P��W;���g�28+p�sZ�e���E,wu�n�"���xqTh�}�;8�bs���5�I1���A�\�칾��|�?���<0��y�dG�?�m���gB�	2H�Atv��9��v��M�	�+<	�J��#��4�ʌ���K#k(��(<���F���(�pb_����Y(�0d4�Y.o^��GJ�֎g��x��䥧e���N*qi�d�>JD>�Y��&�Y���k�y���E�ӡ�+�O��yP�S���A-L��[8�b�x�&��1��Cj*#lX>קa3v���{Q��Wp�0coV��A�G�����.���b�@��9��dJ-VU5v�i��`~+*Tm5��1D�ǉ���|`8c���g�j�I��J���tt�6��o(�� �FP�Q �No���8lE~��IA�I�yJ%�tM�Z���7��;�35y���Io0-�:�B^�}Le])bK�3��Wx���|�2���3����*��.ĥ��H�o��a�iU� �����eQH����7��0B<v��f"k��*����1���6��~��%Qް�a{�f�����{�w�:�kn�%Yu������2��M���ImF��g�(�JF<������M?�ѿFǕ+�nIћ�L��b']���P��}b*]��+��9� �gfu�=zE��L����s��e}���B^lqgɾ�~S���E9�waTt��/�3n3'.e�e	5�:�P��n�w��f���mB^l��DJ��UkP5k�ԛ�((����6�_h5ع�lD���4'A��(% �#�(Tr�;���8LV���yj�Q�+��е�J$�,�f�#��_p�|"7��#f�G,
3���%Rz38<��B��?�/O�N�����c�sC��x��n!B_!2����~	�~�lC®�B�ɏ�ic둭 �3|$ !��L�9��U;�D{Xq[���u9�ܦF�OV���#{G��ʴ��}O�sT�$g� [#�!�"�B|o���"����a�l���1OJD�'��5�d	)�''�DS�^U̝�=���tH=D��(�\���D(�����"^29K�'���vC���w�M�)(I�%�S�'�� �ǝ�Z�����/�df��B���G����D�`�#��`x:��eT�a��%X�"?ʚ��]m��=�CG4���y![���]�D�<J�!"p���r��iah �E�1�:� e�?L+���|r��	 �q�Nv�|�z�ҳ~'RZS�cw8�kq��T��{+��LY��8jH� �+/����#&\ʹ�r]P#���썐�o��b���,�_����b�Q ��BzGHD.�z�����_��o�o�!ܹ�lHaj!�A+*�]�<�iL��7��G38�O�m?Yw{�!l�҈�U9�G6���g0�$�	7��w�k-���Z�_Qy�N��h[V�uU����zp�� U��Ҏ��J�R��gۮ�ʝ�]�R��/I>��T'V��h����!Ѐ5Y ��{���Ԥ<�;�K3|	��Ɇ�7�X�zO������X�F��@�R��k"�m"�o�GA����j������(岳.����/�4j�g{˫xއ�l���8��?�!`���s�3�����o������(4�8�|i8w)>x�)b@%w��BL/y�|�ᕝ��q �améT�T�FW� ��C+�`tH�q���ٛd�uy+FH�<�V��R��*�O��Ҳ�����C�6o����v9z��·[��`�hq��H&s��X� ��y��(+	X���������}&�֘eh����C���A���f�a(ƻy,��]����	*�P�9s<�W���,q��X��B-�9��=���i�v���tP�iF��BJ����
�Yp7V�yl���xio����-�=�/O��G�"2i�Jq�h�!���RZ-�z}$�%0	���Z� q6G�RA��8�I�1�w�mN� �E}_ӪR@p�%L$��+�Æ���ڸ b���x����F�4
��D+�\t�)\CS��7��\�t?Ŕ�>��̨��)t:����|��]<=�Dk:���5���c�CUK�(#$~pM��L�og�T�`�u��pp�����������+a�'�`{ґ�i��Kw�������
a�u����C��^H�"o�iN�!/��f�A�Go�\���D���o�����7+7�*����(��hA�ځ���
��_�7��ƌ5�]�FKC0vc��oh���,xTJj�.f�Q�HJ}vv��@u 6��u��<rU��:�㔟w��a
�O�{�������n.�a��?���EY�X�)�_���ݦ�/1��0�H[>\�]X�[$���4`��@���G��D�`mAJ[��  ��ō�� ��s�\mKM�"~ �6)JqR�gw/ �1�t:�$qW\�(jS�7���\Ec��}���F8�Wl�B��A��˹3Rt�&uK,�X�e�7�'&<0;�����G�q�l���R\��WC ��IQ�D�z�lB���9SLP���GC���CA�����=P1�v�x�@��s9`@A�)ge�UB},I��Fnf�M�p����H�=��e��[K��j����'�
���NFbsbX�;�����>+p�H���a�^�V�6��*�֭?Q�-M�Rpڹ��: y�Yt��]�g7<�ǎ�`u�s\k_�"�Z aj�=� ���x�%��}����Z��}
��e���S#|�u���'�T�u��REs�j����}������i�Y
��6�uH������A̦fv�� !y�ĤD<���X�)�"h�ԡe��8X��\�}j.�<�]�	ZP�iZ�z��l�\^VUI�U��*vT�}u0���
c�+6����M`�Q���S�<��ys��� �{i:���OXJ}�L�^7L������5�t�%��JC�˝�UbT�Ir�x} �����d��^s�*g��
N���bb����/J���ʬ�M��̢����L���ӵ�q����Zi�^��q�j��N�-P��GB9�7�H��8��&g������I�[�z�	������1��	�os�*m����s/�QVW��S�A^h=�`�z��jy06�z�vI�"���Y�*�7}�ݽ;w�18) J��D,(�r;��Ğ1�����Ue���$bd��[z�`"YBP􌊻EW�*��ehft��K��x \�SUa� �+PR.�!�W�z���3�_U5�l��Z4L�W�$0@�S�{8���ʛ���|��V7�2��(r�T�5UUޏ�u�Q�E�nϲ�?Bk�\�&?hȞ1}5kO�UU�V.�N��"o����
�i�1�$�+���A�W��"$�yьe�ᆶaE�[0�m�B���d�l)f�@���ї��qz�ѢϼR����տ�Ŷr�Z���fV�L>��+�����HB 
t,J*d��}����k��)�Lug�جy��,����*̃� }N�V�H]ͷ+��)v{L��P<��/\\���	�Y�}��f3���z�K�=ڏ�i��Ӽ�:�e��̍�9����,�E%C�8F�l^e@}�h�~�`"0m���������u=Y�j����7�����bT��h�L���e�Dg����_������b}����q�[йm������3[Ǽ��=������Mg0�I�h<K���cJɳF�"y�U;A���0^�Ū�o1N]X{�@�J�)�԰"ˬp\8я���a7��.+ ^�d<%��0ڥ}�/�7�X8���~h��є}ے�&X�ʳ�5H��ʓ���yH����dt�vj+���p�P#s䚊�
���$���pk<���B
`M1�	�OuoA��E��/�R���l�f2V&�� 1�a�{q&��aS�4}"}�ˏ���Z5|#WT��iP���}nmD.�����U����,���`,�Dh�G����撁 j�C� �����^y������%��j���:A�FF���T{Pv�:��;k�����՘�h���%�u�T���9%�����X�D��:&0��DV��̱fY��Q���s1��B%�}&M�/��K�|���U��.�醢z�%�T����=�@섢���(�'����*�;�d��Z��U����b� ����<a�ےG�8��L��h򖳍u:�x� ~�N$Ϙ6��n�+L@�w�D�'8 ZE�l�\��F��8)�D9�17����0���PG�V�}Cn�:�u��J}�S(�~I;M듗���n�'����h���jTq���N�I��'++��� �QK�;�7^��%>{��Yh��))VK.�q��[�&Ǖ�ï�].%d���"�������������Iz*����J���&��}��E����.z�T$��ıۨM_�;���o����D(���	��L�;�%�.��V�2�P���)f����)\?�D�	-{8��2�I�)Cں녓j����gPe�È�0����zv����?���b5-e,i�N[�J�E�W (=�7�o�E Oz�g�_���-�����}������j���B��J���+�P�+#���K�(V�-rs��{D$�7�}��Hm$?�2W��z����rEg�ɶ!�J{��Sc'�3S�$z�z�jO*�7�X�(�M�\G���4�.��Xnncy�^�S�y�����9�Á&;
����틇ZD	�F���~�0�7U��3�l�j�𷏇7�-xRlv�a�����% ���"ѝ=�Irr� ���67�X���\|���?TEV�Z�-#�O2��Po��8!��Z�r2Dz�Љk;��_��N��T���9:���7D�ľ�
Nw�P�w�����6/����k6G��Tм�~X���-����V=Z��sSk�E�3�{$�^�����C��XUV�yQDcm��N{O!��ƧK �+�����&r�*dt`0��nޜ\��#5��싼WT� ꊤ+��ף�}rӿZk�J��&��j显��"8��\�a���]��f���3R��a�:&6��q�?uZ����+g�IM����<����5�-Y$3�g�T$���2�5</z��L��*��CY�a?y��2#	(W[=�|���hT���q61��	���Ʊ��މ60������a��в(��ۗ8���if���gT�A��ˊ�Ԛ8�da4HcM�����m�7�ʭ���;���d�'� a�"�Dx9?D��B���yL������V�� �`����u�)��O[�Rv�
1yɴ�F�b�ZVD5���7��\
DGF��QL+��Y����φ��w��A����B
�0n��Jh�<����Z��$��;1��<c��O�S*72������i����ʹj{���a��<gV�A�j��&Ґ�Cn�t�z��Yu>���O��k:p�G�e��	10��J�9����a���4�c��j?P&Bc%1���!��/^�%�;S�u�Y�*��r�4=�K�;z��	�� _b�;|~8�zI ����. i����65��#������z�?d�Ԇ�1��7��l�Ax�$(��LO׌c��Ds��1��Ӽ�C��s�~�1:��jjf.�������+�4��%�����E����G�)|9������d�U������*��/������N����ʽ�ƨQ��%K��OوN��
I�\�'/0�+�I{��;�W��퍴R��o6��64&D�����2���z����~zX8Q��3f��a.ۉ</΄��D<��uUJ���O��
���q ���$Cڥ�*y����?�H�s�}�AX��6�O.���8��$[?�c��r(i��|O���ʯ�G�ςG����H1�^�"/Kx<�
�\��V�tW�å�0c��гv���~�)O������y@w�=�ӼPP��~d��P��f��x������XUO\�����x�o-�Xz�l���@�4�P���*͵��H��� �����=LЂ�l���ɟ1��PR����`�t���Jz�<�:���F�EeN�S��.��^�.w�HW���hI�]��Y�mf^�+���`l�^�fE� .DB�v�;�8A���)q-��I��N����~U��vA��c�c�o@�{e�H{g����޳6�'����@E�۽T?�gz��l���l�+���§ʢ�#,�F	JUp�����\o�$0�b�t�U�G��ܯ@�T�*� C�:P�iy�#uִX�(�2���9(m�����I��MW$юVޡ@��M�BߊVP�t�r}E��,���̬\'��=�`}���f�#1.���$��i|GY�I��p;���TD�(���D�D�m�U���"8�R�)���z�ݔ/qŞ��k�B%�u�S�ݢĩ�����zJ�$|~Ӕ��8�:�L[��1P�x]�c�^�������i��✱u�Y�N�/a&�T:`K�+��?��N���4!�"�����Fԃ�;�?���ce:! G��_z9���Y�(���&�q?���͌"�9_��!�\�`�r�Y'MU	�v���J�?�p����^����m{���/�Z���O�@$"���x/=�}Mފ�^P�G%���-	�Gf1�PQ��q�BRӵ�������`׹�䤉C��!+�gVXsW/���5�<�;U*�ǵۊ��p���i\Y�IӖ4+�}��7���wf����B����k��e�JI�"d��~���Nl�Ug��gc����I���\z9�%{Hɿ�C.�Av��N}:�F��2����GV�~�P��`�/TD�Z��F�#�.�f�p\`Q洒���)ܺY�I��Rc����
!Q�������^Y"�2՗j�߃�Q7O��"�a, ��ej�P�S���I�W�7Un��*�{-����ŋ�_��g2�Z��S)�Z��C�h*-��z�5���(HSm\�Z��:!n�RIH���(]8�A��<B[��<oVox�,����ߨ.�����d�d-buRq�E��!J�3��������q>���陝�ƴv��
���"�{O��Bq��wP����9�_��{��)��}�"��+B�`�8yj3+හQ�I�M79�囫���4�[	����cM��=���a�1S�mK�'3+�H�Ǜ�`�wW�u�دvK�F?�i
s�_�> �m�	;%�7���Ke�5N4��x>=W�0D1�����SЁY)ޢLϘ
��f��a.����t}��gA/���͸XD���5������_����[��<�E�!a��X@�2�ө�\��c2(�-��8/�O�l�Y LP���w!�Ď[��Q�DJG�A�`��/�m]�ۡ��q&��Q4-�\�T��Ǻ^l��ɸE�Ku�o�[%Z�����8�l�ֹv�wFgʌ�Ќu؈���g&��
�� o�e�(}���oÂT����%_�d��/���@Uv�F"}7���Gct�|<[��y�dR֏�xz��0=k�����]M�Wah�u��]![1}���S��t���f�
 %u`�N�Kņݒ$i����p�E=�j�	[�P���!�ɒ�a{��B��c�G>4���=:>!q�"��j͎�J���u<	, �6#�r�d��͡�ȱz�]�� J�u��S���}9�9���g��Ҷ#3F>�~y!>)Y���\����Tx��OAO�rDv|pQ�u/G<� H��:�]�0 ���S8z�|!v��4��3Z�лs�v��\���D"b��
�q��oy^Q�c}�s���_�i��U�8�$����.�ʬ���K�E�NF�P	:{�����*���hsJ�S�o��+Ǖ �-�J��r��&������F�o�u�X�!",*����ˎփ�v�c�7��<���Ef8�Q��Q)��]��-���{@�����G��x[�$�T�M��/t��2k��3�UE��܌�����$i���i���$�Ƅs� �qd��$2�.��^ ���>%�~=��n묌op��8O��[�X����l&���W6	-Z2�I<2ʕ��ݹ���a
8�x����g@ԶI�]�KTd�o"_��5��S�^���&V��I˻��	F�1Ca��X����i���y~ܩ�n�̠^-�<���ەe��KAV�����������Ɠ<�bY�i�'��;F^�[��6{1���j�lQ�W��\�W�t�-�,�T<�a9���~z9��'�R��U;[Tv	�ʼ��]w�j�����(�iFnL61�\T�a&3�!��L��t��1����Mli�t�7x��O�^~>�sf@��h������^,K�vٱƤ6e9�EMkyGk�@��|}u$�@fS_$��4�-���WA��Wj#���]�ُKf��8��s���U��;���= ����JE}KR���/��۟���vϦh.,�d�^c���M�G��I�jH.�a�2�6�fZ9��7i�a���<�d���d�d<)^\6�Wx�x#Fc_�|�?�B�=I]k�I ��$���I�AB������p���|�Iy��$+�8��nք/�n����%�1O<*p�5�vD��t�%�d� �U#��{�N3v�T��=��C�Ж@�Qn#��+0ya��	�*Dw�6��R�6��qOEqG˸�����I���ƪ�%��n�"���*�����?�z;H�)���9���M�P��kLyGu�C�=Ɛ��s�k#�v.���-��I���`�W�uX�o��H��t����6�B���x�fW��{rf��nEu��e+��X 0����+�.�Of��(!|���e�T=<�}m���C��[��E�]���=�3�q�5|�(:.QS_��eQ�x�XhN(�=}_��I���\l[m�(A�l.τDF��q|C��b��=2;01�H��)U��M�|s�����J M�#rv���8b���|��	�1n�#�\Ν�h#Nd���~�>)}tHGJkK�QGB�&��"C��Hڐ�sb�[��&�֏��p�<���� c:�qH�{���Ǳ�>���.>(�纉qyGkl~3<�X���>>�l��m1z����0��-X��`ɔ����b(���9��,�;ٔ�ޕz��@Ѡ��r�oT�~�DF���*�.��U�!��1� �Y�xMOxbL{`oy���]VZ�>9��"�d�i��6͖F�η�Fmǜ/C}����\��$H�wȎ0�M�I��kJ;�d:2`!�_cQ2��u	�B�H�G ?dyq�MW�B��LK"��h�����G��WG�V������Å"�G��'s, ��[+�X@ـ��s}	�1�iڌG��Fb�\[į���9�����خIh����h+x�/�qkU�mɓ\��$0Evw�)��H��s��k�?6�ߩ�im|O�����5b����L���T�>�� #��&���3?���թ�%F��W��zb<��� C|�\�o���t;O`�v��ڠJ`U�ک}�ɢ��PA�_[H�"
����Ť[@מ�'�iއ�#�39[��,�A���D��&}��x�y�K�䏔���G�Y�.��V4�V��g .��eC�p���_,���>��rU�7�^��m�s���^��؅ܑ�Gۍ42qRP-������(��϶��:�/j�����!�ͧ���ay���r/��Ui�-�ĐݟP�`�}Um�lsx�M�w���r+�Ӕ������cVʉ�?����w��!���0����r����5#��y
�4\��Y�}�S��x+��KJ��s�e��V�B�#(���j)4Х����������� Q��iǐ�xc������)=����<4G��ǵ�P����eM�y��u#��$��A�%__�P�sQ~m%P���ը����'���o�4*��H�t����s�~]4�I�;��61���]mv���@j3=��Dx�'5'�9���C<�ҁ���2�y:ry'�Z��=�'�F��M(��,2�V�J�{'��������b�ǼI��9U��2j#ņ�b����p̄��y:͸�4Q��n�@�����f�E`n�e�\A���6^��C���Ŷr>�X�n���h �X
�	�&��KYI<�7�̋+�(���c�$����7��(�\VJ/�H�ȸ�+�c�f��u�V�Ù���յ�l�Z?eiV�����1B[��h _�-F��F������$��T�	:�5�j�7�<$�9�@
��f����W�G=�g��U�*�M=��2zO�5ŉ������� "����,�"�0u8�����͔d4����HVG~t̚dK�va"if�j�V^RpX��nc�G�Z2�A?s�d�34lJ��jZ��Lp��:b�U�����&���A��P_���x��H�a{rN }l���5���A\K��sJ}o�V�pāb�.0D6.\[����t���Ƿ��B	3�����Z��;�Z�+����\')��7��M���(+ɜ�L�E��	KʫЫ�[nhh�S�h�̫�E��	�����w��lJ�>�rǕN��Vϧ����t�2��%�iv��f�t�AAK�D��8��n��l��9��gṧA<���uz�ŉV���{��m��ȣz��H��8��{L/h��������/Wk{?$DF��n��J�C8�mJ� �1�BL�u�� .\�c���ms�a�ȴB*p	��������^.zNb���J�Փ���ˏ�O[y�kU1�[��, 3�t.c���˨��8���쮾�f�l�'ō��H��((!cӓ����޿�\ŎihA`�yi
d�4��h�{:����S�
p�$�'W�\Mg����ٰ��n�X�����׭	qx�\}�0?�����0�8 �Z%>ƭz�?��WPO4�c)���L&�]���I4J����
K��<�bӴnl���[U/Î[��|R�o�M�G���,Ie� ��裼�܏E�L`�KϴE�B���4�x�y��][��x}����UfJGV�V�%5t�T�x�6
�W
*�b+���!=LUJE2*8)�����(+�y���^W��D�ʂ�
���%�i��E��i^̴µ��-BoZdf6�4R4d��@��g�L 
��k�ݷ��������#c�Xb5`D�G&M�I�#��dɥ�fn�E`��&��d�����E�V[�s��G���C��hD�'��{�t���E�P��7'�i[�b�<xm7�����Ij>���J��H���~��_+���%@�� �ʾd�X�¡� ���eKF&Ֆ�l6t������}�~{���j��j�Z@�W��C��z��1+g�h��"�:Q�3��?l9�0��f.4�'5���P�Q9b㉸N,W��`(�qy&��g�b���Ä�cWX�魇}w̦�2Ȝ�eF�&�����Âޭ�YP^�����k�����YU}1��f/�Ϟ]qR�^y�u�n=��~�n��:��%����T��B
��G���Z��e&��Z�/���J�Mx�Y�]�J�	R�-̱��`���Y��Rڇt'T��Y�%�������ʈ�����^�����U���a׼z���=Ty�e1OYf߈2`?{��7��s#QՓ�&��=�}g?.��i&�	���y�f�\�1�`��gAYI~~>�5˲#q��#��8[�d����nν2^�V�X�����i��u8���;�i��Т��[6�8��q����	c� 1?�>�����t�O�z���Xj'�#�)SJ���3��4�Wbb�������4�c��9��2����v��x����b�]F�U$��<ʞ��������/��X�82ڸkQ�櫪�un}�`����nNM\$��i���_O�]IN����x�c��F�H�ub�,5�C<3�F�Y�䐿g��Y�`��t	��� �t�`��+�5�8ij,���w��R�� `,"��p���$V�����CE}�^�i ) ��Gm�`k<��g� 8[)��"�m���
H���{kG�P�L������S�jOd�9��v�_�s�-�I�A��� im�Ԑ;�W�C�a������Q�\{�TZF���j�|��w�%wa��vK�>�Nt��nmr6���Q��Y��O4n�#Ew?��������i�z����`g�]$&(�v�+�t^FO��_-�q"�t ד�i�y5h3(�R���(Kji����]�Ί���OỦ Ҭ4j��P�A��Stj������E[ɏ1��c���&����̌,s�+>��>�t��N�L؎���<���7��^�PHr���z�M�r����Eu_�P{�Ņ�1^_���%���y*r�� /��*etf�M2��Q�v�Es��w0u�U'����zb{:��蒇���я�=,=�ʖ�N���ak{wG�@�Lc	���ݮ�oB�b�~
ֲ�ʝ<5oG���HSBca"|��i�U�X�����ɖ�ΗF� �W�՛;���6�p���
���V��L����̱�ۯ�K�d� �1T0B�ob­���%Ct���S���7�D���ⴑ,j��e��չ�9�q�t&��HS���^R��@�����;�cd=튳I�S����D�x8$T���ԯ�vq��ŮO7���j�0T�)J�N������qZ���23���ѰjW(e�ޟAEI..@_ ���LZmK��6��1_'G����Ж������s\�� �������7�Q� ��r���N��l��xFoa��{J�W�2²�����rg�F��`�dp(b+����t�+Y��".��$t��q1y4�ƨ�e�^�7F��J�h���Ӄ����ZH�rZ6�=��-l�ܡ���n'/�4�~�h"�)��ECÆ��{l��8������G�F������9/�..�Z�' ��Ԯ�b��[p�VOMGX��A���b�B?��ts��GJO��h<���p��/�%ۖV��3_B��	k;�k~����$�=�>F��b_���95�v�~-�FK���(�F!ڦ����D��������&t���<s39�ԑrܝ<�!�F����%nU 㝂�����8'I�P�2�����|��F|��)�2���F�����l�}ԣ��`�Q8��\�b����R9g�nrb�-\��A`�[7�^�b��M��]vkT9O���l�QY9�7p�8��i�Vg5R�(���Q)�"a��)��ݣ���Mc�ɦ��%��[���W�
���GDuX�/���&i��q�C��e�t��XZ-���J�r	�G�t�	��i:Pc��Ry	+aJm�k� X�P��h���X������W$�\$��̎l�y�wZ=�ގU�q�¿o���0z�/�:R@�B[�ٲvA�˨���h��b�t��� :ׁ"~�J�`��ȟt�|T�t�X��vF}�vM*�b(�x�.���
���D�V:�o�XRW�Zi��jFv�G�����".B]��H1��/:a*�)\�B��B5�����d�gN����]V�&�ʷ�"�k�,�%����-;5YN��Xǈa!v�}��]��NQ�{+�$W|K�	�(�G�\��e�K���ݙ��o�sF@_��>���i�a�q����a������@��K�T�ѴtQ/�mʄx+�1�[9��ޮ�p��&�? Q^ˤ�'�%���sW�{�R�{���r9�bq�ʕ�#�ο�V��D-8Υ����Й�?׶G$s�߶~���8hP+F�,)���Æc�`kM!~Aʫ�]C!_Q O~��߽h��NM���G0?����̤c��*D�۶���~���_� ����S�&=ffV����_����s��6(|�A�i0M;��-&F�3��y�J�D�R�KJhtB9&��-VX�4�c��${���,p�b�_��ۿt;'��l�l�j:?���ر��T���lP~vadW�뷗̈�{Łf{�Ƅo+X�C3R��z,{Tt����x�'z$_n�7�9\��G� i�0�$�K�W�[Z�X)x/x��Y�P�E�[����W�8�!aƃ��.s�2�BK8���O���"j���hN��[`�B��e�'x���).�+Q��������ű�&��6A�<��9�`��^�N, ���(ݞd�O���X ����c�� m+�l�DC9R�i��P;gՔ��(Ht%������䴤D�a�V��X^Q�.��ԁ�Y��W�|x��a�Z�*�*	1Џ-��C%�ң�yB�x)���"ya�m�Y�#��)�$��;ePLUDzI::��B�8/����E���I[�H~�;�H���(H��<Ղ|�}LQ����|�.A,^��q���J5��a��v��jD{�+�e(�XC�7w�$�$�p�"��O梜�(x�L6��9���HMq4�d�!���b7ê����p���*��$�æ7W��?�&7YR#�S����G�3��<���@E���c��M�c�rMF�{81��2 �"��A�@���Y���v�	e��&�q���P!��]� j�>&1�m��24	�\eB��e����֙\�~"�;��ֲ;�v��5i��8�X��U&Q06�6R�k.�GHEk�>�%Ieg�NQ��|-�uIA-\�+���J4��v�b3��~��Z`Q��M#����d��rڷ��͐i�0��wI�Vp��.jV	��n���&�����8����r�{����~��I��� ��y�_��!�N����*6\̇�}Ms�ǌy��1�N��V\��W��]LN�:eq�e*�w���X*�xa2����W=��A�;�$'LF�6�W1!���-�)W�(�<�ƞR�}�R
 ��қ����!ٸ���h{�<�DD\(�uE�M�W�|_d�B���O�Z��
���İ�ޡ{�����>��f��Y�0}_�W�m$j�kg�wgʪ�U�1^?%�Jq=�I."R+�bFR���	�p;\WFJV��*Ao@�Ɯ��5/��JAZ|�9��P��ܺ���� `|8��\�����5f�����cdr-ӭ���f��ZGֆ���g&��J�u�,��
9�_ŠU:�(t����s��

pm-|ɦa�B���b<��2J�z��G$�hn,:�|��C�n����;&�i~oxd\Sa>��Mj������X�3�r@P�~�Vl8�/�Xc�ű����A���9����E�:g9(x;VA�O�9�f��|��y�^N�<�S��bq,p�� ̞1��vG��^���a?=0ӂ1,_J�a�3���gG�=s���Ro���n����)�b�3�6�H˳�?X���B͹Ѫ�r���Vw2��� �o݊�A�KtV1�����,PЮcy�tD7���Dp�/ &���g��5�Z�3���
�s>��L�$�~ ج����$,s���0�7zd�U~�z����D\@�j�[�H*5�d|D�~}���k�d���-���Xډ�HEzm6��'k���:W9�cvCX��C��D�U*̎x&����ut��4z��c�++ip�Cr��#h�|��A�j7ƀ'ߠLE���,�ֽn��v_V�P%l3��i�Q�Ld����Y���I%C��u��<#5�ܛ>�́���Y|�ۻ�������⋊)�(�\z��TH�B���*@�t�XPϰ�p_殑@��z���g{|�D��ʊ�l��\tض��P�s�>4��0���
8��zx s��x,�LyW��"�s���=���`)��HȤg��
-��lk��QD=C�v����8J����âw���Wޒĕu@����F�n�8�|����:T�����}���X'O9�9���!zv�� y���t�m��1�	 �F�g. ��[Mw�Tމw�x�6����c�����gK��54���H�բ�(���Ry ��7�I�n;�"�
2L�#�j�_�Dl�(� o�a��5+��e�;ל��ظ0�f�v��?�W,G�Fvb�G�7_��f
�(C` �Xޡ�`�n��}��w�-hՉJ�^�7;���`�sk�1B�]�nbܶ �AsC���!0yJ^���Ls�^a��O5TȤ7�����$C�Qҟ��|�#q�cF����OI��,�i�Ƶ�+��Uw*�^�q76����*�Vn��	��?V���A�I�5|9�r�Mo,�8��"�@⽣R��p����2��?$���(��ͥ/m`P���VS���<-�/����`#����r�_'�1��_4���\��}�l���Pt���]x����I�����?N�| 2��*�|���-�������#,߿wԛU�k��vy�w�ۯ�A���'")��/�|1��T4*(�J̕"����*V���U��3��QKt�ɗ*-h8'�Ɩ����T�,7|U<�7h�|1�nySWh�N��i�gZ�h����\b�Y����(���Ss�4Π&�� g2��(�T�3�v�t���S͆��}v�ј-�N��������l�4���$T�f������\S�!;`x�ML�3��[ٲmw�Թ���	`!��.amU�-C��Eb�K�)��
��S�i���p_`�$A+����f�t�.ͬ�Q>63������w�
I��bl�(8���>��i�xX��lry˙Ke�c����F���6 	�3O.1�����_��^)�˰���-��Q<���wx��{5����G}��l C��w��R8�7�U�����p����%<>ol�AAi�9Iw�O�ɿu]3d4��0��_���v�j z��yڊ�-u�m���?z�5R�1#f;�7g4�j��ެ�.�ߊ���!�æv"�@�p<�|�o��4�9��՘�'�do�Z�(��Jb���uoBʼ)���)�q�w������%:ӻ+v�f�A�ǈ��@g�=G��Ɇ�����uVʞ�<��.~�Il}���Z
<ybf�<���Y��芯G���<#��;��	�:]��
b�`�=%1���;�R+�L����͂���*I�)�:l}'��aq�A�Ϩ*��c�#�|Q�v�X����Ë����v���&F�m��r�^�Q��K7RU�bc�*U����#R�z�!Gy��P�?���1��i�wP�FAG^�@� 
�Eں��6޷� ��z��Qj�v,?t�ѩb���	���A��˒��`�|���V2��P7&�j]�AXil=���j��@��'3�@z�~G%��N�~��D�y����#����z,�� 	���=�T�?���y�|\X��BdE�0�pz���πۥ��P`oo�*�z1��$��]WW�,Q���!~#�S��LR䰀:�>f�NV^t
�od����&��#_]�/�v�[��k���F�Y����u��Q��t���k���)�y�A��C��Y�+�I{��3~�q	���zý��v㋤��^���;�����+��}z�Hx�y���a��֟~�~�	
��7y�GT3�ȗ�;�P�����Lj��;�/�`۔Q�U��=m#�u���IC�����uL~47j����7�jh�߯�yI�
^�#�t>��dz��aۜ�Z�5N�eK7$���C	FK�u�_����t$>F��z�@YJ	�p?�V�[]MQ6�K4��M�M�b��s��\���7�E|��y��p��7jH&��q��x6����\��R)&�w�B��k�YPj���vҫ��Ϥ��$�$=�����&��5�&�hN�\���Uhw�xS74�����i����,�"4���%䷃�;Al���g�3��f�0�e'�E��c`X!�;ad���),��@|&4^%������%��b���k��9�6
��X���Aǟq�|��sE�����Aq{�R$,�� ��6�|^�y#��G��x�����e���M�J�/�k�j�<Ou2�P<Z��F�B�Wա�ٸ{?%�F����ѬBz��I'</���n@��w⬺nݮ����sl`��*�Dɖ�d��<���K��,�o\��v�LR�7�����Y�RT�m���`��`̝q�ԛ�$)���ؔ��[\sL��T�,�>��il6�~���$E﾿ٯ��Hj�ڰv�}Z	��I4�Ha��M�	��S�HH�*�]�֤Ȯm���n&�h�*H�~3�
u��@ 2M��`�$a�jE������sj(HL=�/̲HF"�(�ȁ��[��v�~Β�t�L��F*<���6��S�6��\,|��[O�;�g���TM��Y��҉$�a"΄3���#3��ӷ������o?LuViٙ�����_�*��4=~컮��k��74R�B�[~-��f]7�Ví|��\r�
2v�[����>�Wɬ
{͏���p�Iٱ� ~Я��쿠����3��z%w����Ox��"G�27� ����@��|����1;bY!?���I)s-�]���q�jfƹ.<U*�K=���tv 
�!�$N�ܰ�Z��r���=���	q�F�)u��ª��ۿ\�N� r��S�1Y�%J�?���Z��y�Ea�]��z��®O�\O���pG���g���u8���[["��D�P��7�&j�/}���ϱ+'�~�����f$�'ک7���w�>�|�`���T��%gu-�p��b��G��V�vC��;�3��g��%OC�-��D�A�����`!E,��]���~���]�}���>-�
�Z�Y��W8S�[��u-��b����?s�"�덮�R�bx�X�1\���G�[�������cD��l�4���y/w7s*��>����-���|?ƺ6��'�z�Z(Me�� ���mv��wg�'D�/4��|Uj&���ԗ��f�@{�߉�P��ޕ�)"y�SU)�)�b�/r.l����yȰB7i�B�hO�
���]00xv��8��������h�D�}�*c�������>d��
�xԩ�ӔD�O��W;�Kh�8�5��pX��G��_�%�sJ:�](���2g��S��i�t�܊���r�A�j�$7��;q̡7:�i�w��7��Œ�7�Ņ�E:�X�N%���mlIR� ���*�I)b|q��Ȥ�@���yn�I��Z�i݂��K�l�.�P��U�T��i|� ۛ�2����wܛ�U1J=cr������s���/%��l�[�iN!?��^Ul*#��*�$_��Wv3���[`�ܻ�J������!�L���>u6�)��6D��YV�3D0�Q��W���9�A�EH�b��t؊��P�R�ng��S;/��ja�թkQ-��yE�ȣQ��ߚ��͖$�w2�'���b��6ƯHy��&�up�����w��rZ�r�U#8Ԝ��V�b�E)�3�28�f�#D
�;8�y�n��rS���q�;>�S?�i�~�H�E0Cd�}����{�^'�.[ʹzyѢsZ����X�^�<h����!ԕ�t��iS�֟��P���T�S�K��P���;�ѿ����]g������t�-DMM��QA��+��h��!2 �;�WJn4c1��<�!"�]�k��5��o#xj���L%����]`y�� "�D?_u�~)�����M�a����Sd��%��5�.u��L�V�͊*��KYf���{s�:N>�p�����<��"���P���̥vi�\���Ks�%SO4F�����#��H��XB�5]|p����؅��>4RM�ydꬦ 	�}2@7^KC�+�o��� gվ(T���>��|;�/�F�uYCˬ�Z�H\wM�V���kq�ۅftQ�(B�����tb��.2՝Ң��?���]Xm�o�@�����&�Kۊ�����)ɀ��o|�{�����cIrv���}���d��5��������@L�[����},	�8T�@���a�zp?x�;v[�ve�7�xW��~����[��#�>$~��s���h2�J������E���� ����"tC�=�o�^FYt5���@/DL�wmy��S��[e�`�,f�֗�H��lt6�)X���v9�8<�_8S|b��fMwH����'O�+|L)P{��><q~6��lO��ܼ�^�dl8-��58=��o�}��=���pV��,�4j���a�ܨ����;�T��[ؖ�bE2�8��H{�{�4��K1p4���8D��o��U�;�P~~ڶjˌ�5ݯ'>�U�6[�E%����p�z\��ZF�2}�M��eP��*i`ljHB�m׿�<"ACzr^�%%���Kbi���N^�xm_�q��f���Z��)k����S���!�K����u��P��W_�r��g�`r�\`�TrQ���w�]�E�K����\��1�N���zb��j��dB��a�f0��ѽP�ͿC�[��-挈�|<6��nI�6�PJ����V��5���l�a!Uyr�t�fqHՉx5�s���}�5��e���gɊ���Y	j����I���<�v���C{��C-�a#�C�[@�X�~�D�j#��ͺ�$ͻ�n8�S���cq Ih�sN�D�>u��Q����Ng�p�k	Ƈ�xF����Vb@W�T�[���
� �p�u}��ӭ�|ub���UZ�H���x g|_�4:�3䖪\��WH��@�^�U>���9��{�:.����Um;U�w�b��{�뼋�D9�
��	�p����bƔo�����]X~0�܁�e�:k[��x��O�{Ҫ�1�(�&.1�EK"��1�c��H�����#c^Y�����Z~:Ϲ��X������d4��Ռv �I˱u"y�����1+RW�B>�]�s�wx��i�<;��=��i���;�Ơ��&�焸���]���*o�\FB��[�iM���Mqp��	i�ێ�)�6��kv�������y�������&΂��m��/�5��m�u	��v/J�S���ކ�G����OR��ZØ�-~UҊ`4["�t �N�M�;���]�3�^������1iX��D �#��.!��e]~1�Y���7t.��T>WS���,��3��T�ٺ���uG�8�rHw�75��N@*��GGPٌ�X��"Г����rp�p
a=�8TG�!��R�� �-�=�F�q
u�uC��QE�N�tx7%3ʴA�G���)^´JO/�^�$�9 ��������sI�f��dʩ}��)�?���[�a���9��SY#�>P1�7���9�_�{�[�����ķ���O��\:hS]�I
���Mw���ћA��}>��P�\�X��gz�[��vZ��,���������<���4�FaLm�� ��c62�JI)�󚩹�||��p\%�!B��}U��>���4�N|� �i�܏�C��y{_x>k��~��U�ݰ`���K7�{�(����ZԽ�� �M[h`�m�O`ܨ��~��������>p�O~�K���^���tಓt0Api����-3� ��vpN�\�� (����~mx��}�����Rӝs"�}pTt������p�������.�
�Hy<ٽ?g�3�GR)p��wu�H�v1<	��G�L������%�N3���r��6M�U�H{�����M?\1�;�Qp��	�8����~�8���Q���~��P1>[>%"t[/�k��x?�M�t��ڝP�dIFi�l�`�Oh�/�)�7gԓ��KM�wk��<�[�*�k8���d`�&��!(Aچ��C������~����1u��,Z��� �j�\+JqY��~`9�Ό
c�0��8O������b���M����hlt������%��,]'F�W��[�"��7�2�!1="q�>:�:5@(�eF�ce��{"n��V��{U�P��" =��w ��Q<�͋N~A���鿑�I96QrHAU\^hN&�>1O��C=�|0�e:���Eͦ���>��1�P��1��E&��]���I~�7��{���C��� V�W3,��{O���M�=v�����L��Z��p;_�`��c��w��E��-��u��>�#��]&V�����Bi�\7䤼���$��Om>󧚶ޖ8�mL�2f,�ö:P��|橛�&��!ڵ���	{��b4_�E�_��V�#3�4�l��	�X@?��x����s� Cz�OzTھ��J��������.楏'�H��r)�%�6/{)w�!K{qJF��y����3>�Vb!/�q�I����<��n��f=O��"�ldE~��fT���5/��瓜w<���U�g�N�r��P��PN;r�6/�'���:�P������]�G��A&�r�w�ݟzJ�`<nL;F�*J�U�"l:fY�&�w�ݠ�v_�$B����ol�%#@.�:D5���yaz��u����<'��.m1ƥ!�	��^tv���@���n��EY��]v�5�.��Y�(G{8���Q���Nu=�깭�^9ᙫ����I���������Y�����`P��j��+�w�⏅W"�a�
'0�n+D3����Q������K��t]A�1:�'x�⊇����S�G��<���\�CH��L��m$&u��v����h�����U��h�*8�_�[\wI@�ku�0g�Q�!���;2�p+3!7J�ж���̊JU~����q�eRH�������`X ĕ��]��>�"y�(M�Xv��=�n���w{�)DL����G־ƭ'dat[bƄ�uK�;�S�u\�
�����gY�\�X
��o�d4:Y��Q"�Øf}N���]�%��91B�chCм�M�i}(���.>bW�Y�p��ݢ�Luy�;Q�Pe�{�5�8rK<�
IL��'B*���f�&�j�Q.H�h��]1,^q�<�i�{!0�N�.a�d\�\H��>�Vl�щ8�-�s�� �5�^a�e��~,�^����y���ڳ�E�F����������e��փb���9C!2*�'~V� ��r�i�e��|NA���<���Kb���r�*�w2K�{5�����I�o���ΚY�"F��X��S(�AY�"�T���à4�O�X��>/���;}�>�~s��L��w��S�!�g5��\�d=t��>'����jmCf�M�LZ�_v�^�.|�����̏�pui\�M���-Hw��+C���wI�N:���[����a>�y}��ƌ�͈�������c/ؤ�W�Į/���i�1���	�T�	��=�*&�B���}R�`'�1��(��3����d,�ԓ4]��{
!P,V�EL���!.�c�Џc�c�n�\�D�?-��������'�G�V,b���,Ŧx$j�U�� +�~'�Mp�mD���<��!���Cf��[�a�8;�4H�T��~��������z*>��\#�aAQ`A�i�ډ��/�q�x��?���v�u�N�w7����<�Ɗ�5��ހ�:tX��ƥ��"Ы�U�τܽ�
g���X!+/`|���vdBsyY������F&�������b��wNo��{��W�B�`�{� V�0R=��b)�}��%ĝ��`mD�M��9�R�u���_�����#We��4x�JL��NG�(勇*���&�D�5]M1d!��U�����b�~�#�4΂��w��y��gCֈ���߷����B��+vW����r��4���(�C��.�(5���
Y6aYurˡ4z�W���E��Mb�!*킊o�p�8�_�Ջ�|ߢi����4���%������������P `v��%����<g��a_ '�F�c���ǃn�[��l�!�h�oTk��7���r+R�VM�/9�]�q1�7�H<[+:U��A��0w.B��Ga����I���T���ԗ.c���������zV�[$X��e�*�ײ��D����#�n�)y��Q�u�8��ޕO0��8���!d�1���*Q�y�$�y=�;߈*9�b]g��>�]U�3�;G�����Id&#�{�T��]a�^��)s���4�,�F���%?i��u|�w�1.�����]�\�^~�>Z��Z=D^V����9O�q���i�����g'1Q��oC^����9?n3Dck�!��b0�J[A���]�K�s�!�d$�{��Ɯx��M!�NM�	�����ũ��T��:1Ad��|>�F2=R�R.aY��`%�0�;C&X���㵩X$tm�E��ǃII�|�M�~#��2�}m��rM�NrX�XG��;^�,h��A�G�C��`
������j��cN�HέRad@Q�F&d��o"� q��s�Gtl�riû��`�r�5�����=VڽR7���CH �Y�"�2�k隐y��ЎSV;�g߾��1Q�4#�����Z+ۢè�Tk�D|f1��� v��^�:=@��jXݣ�@��@�0e+�� �y���]��
mE��+|�ʞ��`o�h�mw��w�?{�$���R�a�����J�mw��vS�^�SSo�@�^"���K'�Ȝ�v�i���?�K���9�TJ3Wg�f�g�2�M�ԪSFE��_M�Jy���^V-���w��v��x/��\��
%y�W���
�_'W�-wxzΟɩ/ζ2H����d�k
��w�N�t�#��'D��z��/���`��/���=��c�
��߅�2�.@��R����L��2*�u
�رfc`:�����(b�&^?&�_�?��qΐb��.�p�B�4�&���>�����G��UG�4���~�X$������"��v��o��bsÜ���+7v�Pt�\�ȷ!3�]�`����s<���
������*��� ���;���i����`��nVXI%N�t�RQ��NBVG@�Q��������������L;]��\춄�RQ�єOa��%N�۫4�z�{��3� |B�����.<��ۈ�i6�o��tEC׳T0sS���*��}��U�Vq_>nW��gqcp�\$9�=Nj>�� 8"|åW�h�-�*��A�f����*�`�ۧ�?�*�ά��C7	'e��&��*�4���t���S�S}�����V�taTa�.�C��?L}�v�"�z��s�n��SCs?Ű^UI��\�sH^`��Kd܆�wXV ����}��h5��������:?�n6�T&��MQ^�ג"M��c5	�q�Q��8^4}�̈́��}��r_D1���ѐ!ZQ�ٱ�p�b,F�iH�j�(���r��r�TB)����۹N3�)���6B�i\?��e{�B�aƸ?�2�3z])	@_�UH��cX�A�2�Y�Y<���C��f�r({72Ef��>zl7�ŲD�;@e�R��>X �ߓ��RHt;ake�������-�J38�^GIT�*κi{�߄xђ {HC. S��w"�^x��3�÷���8ަ͎�|�^�.ЋAiV��!k�Y��dI���17��pe� V]��&�#��77R@
�U7�UM(�,�S�qn���LH��[ctp�	W��%�Ē�ׄ_v�TG�tJ.�=7ص���5��l���7%�����K��$&��/�/���N"��lcc��;��mn����VZW$Wit��ZA�/?����M�N���M,(��J�kg5����,%$�Ҏ�=#���}�1��W���2-b�ɞ��Q�O��<\��wfɒ�4�㤊���_��7[�} t�:%x3�6�԰`��ar��U��XF�\�*�q�S�_�E|��Z1�����Pq���V���1����Iĸ���F�\��k%����x�Y��3Q#�@pg[��\���A����b������[�	<�&A*���y�����;�j��$�ơ��5�7���_k�@�#����٪�������?A�T��#����D1�n�5Þ$/����#���<f;���~�����D� y�kC""��]��- �דd� ��/Z4c��a�I�q��[>�w ���|��ɣ	;?q;��]ǂ���uR�l9U���. C3��S �0�;�8�J0].����!�J�p̐�S����ւ{>r���4�鞕�ZVP�'('#w92 N?uQ�W��2�@{}�/��F+�;��߈W���`̚A\�I]XrN�h�Q�q��3͞�]��U@_h���nV�g��B��#�p;XT�����_N�М��Wٰ
]W�X�=a���r�%���pf<�,1��щ\�vz���_��yS���3%Ɯ>�d$��f�/ k4(	��X�tv,LY�saGy�����˱�s㛓x�:��^GʟqJџ*�_�у�z��V#;���K=}C�籌p1ϊ<���.b~2�
����.�VcD/����
R�P�cb=&^o��?�n�S�1���#���I1[E^��1� �|���<��1���� �Ɋ������Cs�d�<��K���aa����,B�)'%h

;?D��&6��'V����2
ZN7�T;?/�72ぇ����'	�}TbE�}q(��ޱ�+H?�"�����wl�Vsw�D�@
��yR�������,��o����;�j�����
M�nu��ne)&6��2���.��`g�9�H����f;�C�=5jBբ����JW&=1�M��Z3N����r],Z/I��0�G��z�$�q'�`m�$?�/�->�]�|f�~�c�\�fO��:�\��_�dKX`�7�����U�_r>�C��_��O���TfowA���T�i�A���i��>\�6��c�-~�2G�̑l7g
�&-T�J�v[�Ю/2�/�2��"���*w�4zd�g:y���,_ l\n��A���t���m���=�����B*;��%?���X����֖Ú�X�5�j5�����n��(������oIr�|����F4]�,Ў[4'��nRWs�����Gf�e���P��fĖ19�� IG\1�G�j�^m��y�ZD#}� ��{-#K'
��	��7��k�|�%�@���d�z��c��b���SG)�ث�?�t��>�+�"-��Z#�Z�M�Orݍ铉��.��ݚKHd�%���J�������-o/䅕>D��G�vG$�s�Dw_���7A��HV��*��hFu���dg?'^��V*��	�[���c�2~���I�h�c�.m�Q�� �~c�(�rx��`Ο,T5��}��t�y�1�!!x	տ�ɯ%���\G�KJgR�`��G�L<���ӃZ����2�Qؓ�p�������3��`��1X����9o�2��`��x���c�����B��u�qX��(�J�j���Q�@@���pfd5TD��a71���^�Mb���ʷ;�ǳ���}�n����a]'[q��"OE�=�D+7Gx�!��L�]��Q��ʥ�{���|d���z�vs/d1NUO?�������	�0���vi����M��š���y�!`�JqN'���ȷ@oe���Mc�d��}�[0:p�켸�����bC��Z͗M7���e����pc`P��s�_$�,U-ځ���['�L�M��u��:��6U�e'�]r��f1Z���q��l�8h2��G˄q��>���}�@WE�L�z�C�\���A��D�� 1�����b
��!.D��|"U�����5CV��de��R������P;|�^����\[�(���r�V��B�I�I��	�C�lF�t��_`��K�]? �|��LRnZF^k�������!1R����B��
���'�J~�u�,͡����N��epZ�Ǉ���ܪu���L��QK!7�a�8h�X���Z���m٣F���V������J�ϵȕ�e�iʌ�U/ёM�(�
�}��S16l)�@�p4��o���ȴT��*�7dȎ��o��IWE`������]t!��nd�]��YM-�����e����F�j�2(��=��DI�R:s x�9��\W��8��#�ZW.\�[�����mn���S5�uu�� �`o@�0̚���<(A����q�2�%�Ta���8�K����h���r���w���x6+P܉��o�HX�'\�����nH1�c�&,��Di	��h=�/rc�o;8�ڵ�i��s�aà�TN�\˗&��k�[�=��-_9p��p�m��G�,��"��:n��#.@킢�"/ҫ-`���Q�%B�CY����i��]�	BIc����A_`�r[Fʅ>��Y�K�4�	�����B3J�ӝ+��%��<�>�������_s�6l�K���Fy�k����O��Y���N*���?�=|B���D����L��B���[ڜ�=*�p�!�1�m�QZ�{c@pv�D��`S+Йڧ?:��H�ud�C�nP'j
�z�"`�$�{>3�m+�
u�������S��5w2�mr��ب���s��X��rIm��K�nTS/��e�?$���Z]>�g�x�[����v�6qXŏK������R�$�t��q"%�����Â}x�~9�Vkl�G�����S�5�*6�ş;n!�|V�	U�FQ$ޓ̻�z.ߕ����kEW`����W�;�(�6 �tYhgda�cs>ž_4ۉ��	Uؾ�h�w�W������D#J���Kqh;��s7��ς�TB�_����(�G� �^*�a̻�0]�T����z�$ә��d�c���_�/��W^��Q�tj���Q��Z�3�w!�0�t$�v%yOX����.�h�K��ltg���(H�.&���Fc.�1�U�"ݧ�Òc�� A25��zvN�J6���u��]_��	-���=8���������� ��vk콉u��r���-?��-W���$��.�))��7���8@6���o����ٞ`����/�S�Fl��̵E-xYS�ق&�1ӊiw[�"���_�r�Klf���^�x��h?�.�7Yl_v�'Oz�Q{lj�izюYd0À�ҦY*a�Yz��$s�`���������.ԧE������h00�+��1����B�Lu+
�� �K�e�E�SGnŶ�/ޙN�B����_I�'���^�~����x�t����o��oV��y>�9'﷫����x�����	�+���w:�#���"�)�V���r���^���a�8�((Jw�Y
��;�w���}�b��k�:\(�dc���C��(�9�Rx�D����y����0-P��b�V9<)�q唌���S9�e�)4�I�T[:ߖ5�}P)�ص���M��V����������1)����Hg{�e�q�_ރ�O�Ș�	H��+�`�26@>(o�{Պz��1�|�4~|*��e��E콴Ug�
��IS&�{#�pDG�|�%�B$����l>9�8N�� g��>%��A,����68���;�Pݬ�K�Ԍ�D�V:��O��\^F-��|�֋��R��Ɖp!�oc�=j�y�g�+K���( p�F���l��ɩ54+c,Q�\��s�i�|Y�? ��:۞ÕW��f ��h��٩o�x�a/���HYoW���M��1e�Zlֶ"
�'8�fh���NJL�A��SW�:P��~�������{�%/���j���s2FmS@Z��D����i� ���(�P��s�%g�NN>㓬�@�0���^�9����k�K�e��g[�M�5Ⱥ�/�1�C��a�A;A�4�~�j��%wf��9�����`3G��w��l ���d&���~\�
uٹ����ܠ�?ɽ3�>�^�y�B`/>Z�j~�v��5�>3V�؆Ѝ�wp���a��p���zdP��l.�"�����.$䗵�o��$�D<��x���s9�7��qh�g;��,�:�}ᔦ��&�\�.�%b�7�h�?^g�v�.��8������ɯoz�ݍ��Ds���㛔�����"V�1�S}��C��)ԄD�X\�6�Y��bd�	�2�:���������NbNP��x� �J��w�A?�5�`g&O-�i�'�i��J'7�� ��� ��I�ܺ�<�mFݮ��o$1zw��KOm���\Z�}�y8a'e��  �>��f��҅��g] :���qY~��S�..�=	k�4����Y�QN#���(��Z��-�VtM��-��#f^-���o�	�s�{��pA�t�j&�L����9^�7��[�ܗK�n���BN^����\]b�QM:��.n	Z���}+���&�}\ �Dpq�n���\�$������-������vC��@��z�=���u����5�O��� �H%���bP`ٍ�/��&��P}>�3D�)�㸛P�-�,�//�[���.��o*��M̹=z���r�Z��ٌ@hB�v���ҬWP�`���!����Xpc�zd�D+��ROS<��ZWٻ^"������`�b3&;5�rae-*9��J�ܧ���
�W4� qZCM^B�X�m^��3,�F�ܲrrк�ψ�>h��{ԭ���<#��G�@�%b���	��8���.�v�� �_���9oe(6��0ϰ1!��R?#]ŕdǕf>��4����#�q��^2���4��K��_Q�`�Vo�ZW~�C�H�"���)��9�4�)^:���ք$lY���� S�Ǚ��@����y�'���F�c�{�@$�hŲ�ທ��R!�e<\��R�m�d�t��wkz�h1���S;��Z�sg�1k�8��6�!���d�\���#b\!�\&�e��vi������R�p)�v�!?�*�u��J)�n�2�h?�A�����U9C�G�	]@���6��
z�i!Ԃ$���Y*�S�G�.IOR�̓�}Kl�C׿+"�Zy/��Vv�<5�4?3��W��n���gƠh�0=�F����������;��_�sr��R������ ��:���E7J��D��<��2��3�
�@J��1�v����w�T�9V������02}&�٧%�;��.[Tqf7ƿTV��p�%9��C5�����<9���O|�*����7��r�ԑ�正�NMl}Lھ�tQ�!v�ˬy���{z�<�s�!>%�@�E7�����z:���,�� �Dc��1�w�Y�P�V�����鼷���8Z�,s�"ݕlև�)^��G���U
R#t������(�w�������e��a�E��lD�>r��1�o��W�y��x�ѕ�b�w�0%�DJ5y���.M.^�s�2fe\}	��B��V�.�I��x=�_����ج36����ҿ��'�J���rT�1�@	�/������A�L��h"���#h�7^�=2Cm�Կ�i�[��˚�5^�#�m�h��e`eA�@'�]꽁}eI���ȸn�v��3�yd�r�-pwm%���""��j{|�$+Q�¥�O��,�c��V�8d�`��tQ�-ƭ�\�/�����칫&��!`R�DX5������g�N�@~�I�>��~�0Š���?�%����!�AP~�@�4���J	���W 5>�;#��� n�nx'����5?i�>3�4�����.$y7Q];��r
v[M� ��բ��E�xTXnʢ?#c�x��L!�3������︼rXM_����՚2�~�w�ɰ0֕�'B��F/��>��LbT�%>�i������*��j,l����z�,bz�F:)��3Y�Н���^��/Zh�oY��h���Sc�6�vW�G۴4"6����^��0��� �h�f�XF�sV-W桙������T����Gk���:jLG@�"�.�7����?�R��妤�-g|�{��_������:�JO� d��Ji[��q
��}&y�� ���T��)2>��]��`����?��t:O�#��p9���ePe޲�h����#��7�G�b�&��E'�+����j�Z�Νec��qvO� �Cy}���t־݋�_�={�1�5�^��~�'�I�@e�|�\�h��2�Ww@4Mlk���w]��c��?�6���Y#?��LӄYJ��bĦj]'�9zN�P�C^�h�>�n�9GX&hNU�}����n�h�k��QҼ��Z/u���_�y�J?L�|�hT�M�����A��c�e��0з��@���ⱘs���W�Vˈ�v�̓rݸI�sH��Y9Q�P<^�".��/�H��U��A82�]���+��P�'h���@�BՎ}�W�޴�<�/f4�iab$������N�R
E�(*v_�8���na���ĸ>4���b[k*��!���Nm73���,�4�j�ͪ��v��KH���w���~���1�|JjCj�<n|�5��YջC�z,>0e'�!V��YD\�SWP#/��v9a
�iŖ�x;T�N�(�c�9�19�~�&U�����
�������X���D"$�f.L�F$գ�Gv�ѳ�U��+����]���}�h��D�����y1� T5�r�?���j����;6�@�\[g��_T|A� &��M�p�s����א��Kg�?Cz��M��ɻ�ڿk���w���c͖ɚ߱�O%�n'3�g��6k�>U�����XD'�\�Kfo]�}#�M.Ｆ�\�ί�_ř?�c���m+�LЌ��I=ђs=�|��
�s*�h��c5��{�d\D�@����/�P#���e�s9B88D7�a�Y��;�ދ��o�.;;� S�~N��5)�e�3���}�'C#�v�����y f�Suk�\�]��
[�"Wx���t_�S#xV�� ����S��j|����0��O-�A-*�A�]l]"N>~�>�[�U�9����[��֖��h��,��c��E�|��e��2��D{dMb�P*�gk��,F���p^�>ͨB�8��N[F�wݠ��v\�O�K�D%2)pi���;���5���D�ֽCy:�w5��t�g�����g��=/q~` D��C�H�l�j�-nb�~`3|<�)�Uf��U�ܪ���q�U9��ۂu-ۣ7Y�M�0�� @U�z!(eS��ህ��ۺ.�abGF������6i��["��^��B�G�
f8=h�l
�Do��N�ǲg$5��{�T��q���?���D2���TC�*]$�}"�S\a�S��SqԀT�"|�n�]!�����nb�[0�D*	MTdʵ�O��`����E�����]V[�	J�;��3�U�y	_�%2��2
cc:A=;�IG��)*�s������\C����L% �KxF�`$�T!3�[�+mn�'�M��?�y2�4�0���W"� #�M����jJ�*�p��lhx�?$b=.�ŗ�X&3�V�rGh�@J��<�p7��u���o��7�����D�[�6��+L�?U�i<U+&y��0`��k��r!�X(������a�&��&���ع��K�B�щ;ƿQo�%�O��z1�V|H�	vq�*�k�AU�� nG���8���y������qgL�=Q4!1S�v�_�&@��ȵe.
��8���;�uM�qۙ�n��Z@:�]~q9_GiͶX�-�2ʬ��q_���g��X�YƵ� V!�X�.hБ��s��!�YVd��� �,���q{�i��l���{�B�Zf��*A��� ~���`4��)A)Yj�A(���ʔշ~����*w�R��ڜ�c���1%����$R)K���"B��[�F3F�������E���]h}h@.��+����xB9 �IB4�K��8���t0�
����$8aa���1L]����t5�ā�ᢩS3�+-Ż�P&�;�G�(V6��~�=�pұ�Q	Sj>n�
������]uhl����`2��n���b~�i~�M��{�Q��G��`k�?�Y�﷬�H`�>~��4��.$2��^/Ы��22��즚�N�H$��I��Ć�9�q���}��i��-�D5��ŵ�������9՘6��l��q���j��{Z�i�B����E��r{���&�s+��'\�h{�d�x�uW8�� �`��О���a�����w��ˣ������#x(��7�.�{`�m�H��k8s�/�-W��xil�K��s�Lw#�ho+_�4���M��ƌV%q�Q���]q�!�k���@r�F���{̙�Yog,u3D�u[n�rx�ʚͫQǉ��:�`Iْ���Z�%�	�<kI`��,`�̀	���Q��	~C��>��,F��m?��d���	F˵D(��_lc�w��.�Kp3��*(\0�iG��P�V��Gug�� �"���͜͞�(�&�q�+% $u�6�"�/���������xD����`��S��uM���b��i:��^�1�2G����������nᬸ-�:�a���J���������H�xK7f�<=�&3�V>b�����3�1F���~w���'p�:�m/�o7����v9c��\� #|��뎂��f&(���<���II����/)�a�/;U�7~�I���)~�Gx�ZAsU����n�h,��r���	d�n�y��liGr���X���(�ՆZ�^t
x�0����/�I6���qy&�#w/Y�R)袏�v$aWF�,/�ns���j-SW5�d�g�?��y��D�5e>����g,=��N�ok�DA&�,^� G�s�暝*�LhXwP�?=�ʒv��^&��r~�F�I�� ��k�y �+҇��9kFx�wq`���[K{��(~����xn�����Ekܼ_1����u�&�i�>�Oy	�{.a��sI���b����[KOo���y¦��@~AF�2�53=�b�vQ��=AHE
?!��)d&��hG��W��1$�Y	=��l��b5�u,��8�v�d{���@s��	�lZQMM�� �ݰ�&�7��wH��{��i�1�g��xB%�Q���C}t �̊bY�D1p���ջ�-��V~�� �-�
��k+���:�xJ�kr�	�Ym߱6ϳz�oN��b�\p6ھ�s�r��P��M���O�7�~��������%����Tc�2\��K�׋�	���!	[�c�;bv�J��D��1{�75���k�x�1����|���y��G����Q2�]�e�Z۴K�n�;,-����}�̘��H�O��W��ȩ�0�bi'���O��\�]��ڼ���nt�7R�e�>�+��ak�k��#����	�|m$ܣ��ͧ�F'�+��.ۯ���Xǅ	_[�r!����qa�o�v���<�új%�]o�mEn�؉�D�f�cs��>�����9?/r�`%f�ٺ|6��@ϼ�A��Yq�?o�E���@�k�w�[#=�n�}��>��A.�����q��>�Ƨ���NE_��&S�16�08U�����V��vi��]� �,�PT�`��1�M��dM�QD& ��ŨY'z]o�p�V�1�"�=%����+��ܰ��D���z22�[���yc��]D�|�x����J6e}�՞'�Bm��Y���|��~]#�o��O�Ѓ�>�����_�L&v�"bA�$��A
 �(�ͅ�����M���/.����n	L�v�:Bc*e	���y:�|q��ܙ��'��R�&��⨇�"�*��e�P�1#fӧLh9Q�lzrW)hȩG�!_�A;K�K���A�+9;�)
��=r���`8"���0/�`��Mj�0��2lv�۵�q&w�� �Vzt����z�/�ux){O���L�d� �O�S�$���!(��t�����\�E��{+�CʛQnO� �=��?ڨ�
A��-S'��>���s�e��&NM7��UH�m�����UZ�U�� �Cpq�_)j���NO��/?�"�t�ԍ�W�-��P.峗Myl+z�Ƣ~�ҕ�{��1��J��X�ㄴ�٩�n1c�r"#������ˊ�A0�
�~໻���r�� ��#�HM�tK��j\=�,�ɾ���A�m�-���z������������R�a�e�B��'8D�՘��\sf���ӖQ���t������_��ڪi]���`ݴY't����b��Gk#��Q�\]�Nʭ4Vr�q��P�שj��6V��P+Fׯg����b���T� �[��{�߻�)!n.��ق���0���Ŵ�7*���~��D�]ٜ�i�+8P(�'xAK�]W�̫�W?�����?g�=�W�3�v�S�l��vX��@9��ht'u6��z���H�S��/���H@���$��Z$�򏈆�Fqw-2��˻�k�N�JX h@��/"0�_t[����#I�L�A����7F�]�~�I��""�垩��ؽ�7E���q�k����T?@T����6�Rb0���Ӊ�ef����R�]��'X��Ek!����I��D4y��GZ/y��0�_���L���
���L|�9jG����vaCږMKa��@Y3Z�"����[`���\��d�|=eͤ6+G�-����3���R�"���4D�pl8ώ���1���z�w��j�hb��4�e9Y��H�1����t9M.�Y[q�A�p;�!;�2�&�I�X8,�#��`\��AM���GX��툀�8�Y��Y�x�NCQ��C�m��*��F��_ȹc����
~����k��,F��ܱȁԣ�V�BCf��R�-w�a��g�4V��`��6�x΅	V.*��V@7��Zt-V�q���z���K*L��^����*�� �����I7#pv�������2i��3t�d�~p�Ԋ�=�k֮<�²ֱe��K큫J�޿+�F��&ج�al9b#�k*<�Tz�K\!��%�����	w;�o��u8L�퐯$X.�+�sI��<7-ő�\�z�O��TAɰ��::6��BT�5�(`�EOg���5飸+�J�-��Ti�ֳe. a �,!T�
Z�gE:Lg���y��8+�KN'�9(��1O��
�C^lj/�<�b�����Jp�vy��?��A��)�P$,�Rj��ɜI�'�]�q��f<�8����B���*�8_:T���.>�Y4D:��)u����;�XaH���X�a&��_��	�a��$�������Z�	Z�^U!�">�>�p�H�
;����i�s${JC��5ce`=L%�������h����	ɥ���@G<��Y%4W�ʙ���lϊ��萿?`���]]\>p��f@b�Z+d�<V��QI��8Q�f�=d��3,�u;91�i�J��ܠd�5U37�oic�q�[\Y����J,2�(�����e0��gr�s��o�X��k�>���]b��(_¡O��F��oDJ�ҏw�7H�5A�i�,�'�D�V���O� ��w�N��KK�9K��z�8A3O���W<��cz�<��(�)~~L{�1V�E@�ߓ���8��JM|���ah�@�o�ԯj��5�)gB�C�w��������Y��-�R�ڗ<�A��a$~��jd�D�������[W-�	(��~��������P�0� �gGV
@fY9�����oo�(mā���g"Ÿ5h�v=��)8��P���j��Qt�qZ�P���7&c_��!�*�gLߏAN�v�$��R�e
`��7^Ήv,��\�鳔f� 8D���Y�)D,+Yǁ�.�A	QdPs��Ӱ���	����{L�o�"�=a��-F�O�G��e��%%}%�^�M٧$�( �<�&�>�C����li�^�uߘ�T~�+��S`�yC��%p���eNk���������T!)(C�D�7���^6n��1 ��Ҧ K=_͜!��C�>1g1U�C�O��Y�ޤ�C¹��Q�O�,��i��"��V0���A)LU��,&`��*�~�ߠx\CHZ	��r�o>�r,�d�n���j��GΟ�a|隙��i��/��Ȏ��Y7YR-i�:�=�%I*<q�������^�ߪ@�kx���`�}�C8ٖ�k(U|�$�C#�d\����TFr�,�}5O��W�42�>�����lϋ��P�R�v)2�1���#rd�	����tgH�͋N�O}\.(�����n?���&du���X_�hv�c�^)^�?f���9�]Ha$����6	���7���I���5��l1��!F
_��٤�^�;��2�����~���MJ���Sv�c*�r>v�Z~����i��t��ǚ�;��~|]�?7m<z�+�+�;��2�O���#���άO=�Q��]7t��F�e���(�3+ kIP-���V��Gi�P������No͈߭�iҲb\3�ͭ�;MTCj	-jGѐ̭��%<ᝓ�,�sH	U�OӖ�_��@̔B=Ӂ��R�Kp�K_ݽ�dwdc��SQ��%�wh 3�y,b��s��M'��}����f$�+E���6(��N��m��3V�h�	��h�vN�����?N�����n��#��ѡ��� C
6�ֺ�2�'���(�B{L�۵���v�l�OZ�G�	�Ӽ�&g��a܏�4!�i��DvL��F�ݒ�F���м%U
n2O� z��*/�}����|
��[롋ʟ��E����RӜ� z�;Q���!���O� |?��[exf�
Iw��ߓВ#�簈�c;�ԡ�pe�elt%�h2`�E/:�����S������[��Ͷ:�B��=����G,�ĥ�A%e5�l�:�j�x��)����e혐�Y�;nu{?P������ҝ��,ӖY��Q�r;�o�f��K���g�1���k�|}���]�Y0"Z��z`@{�h�2��zD�L��w������aw�ޚvq���L@]z���#�f6�����2I+�'my��z��������6�Ӕr�o�L�'_<�SezSd��ѩAӞ��c�W�q�ط�i��l.��n������&��81�K��N���&b���ج��s�WH��ҳdZ��1��T�f��M�f�X�xBxk5ٔɜ>z����7љ����v�mZ�����3k��*U)�W���.�࿘K���v��|�n<�)����e.����5�WW�����u�-[����w�p�}�a4���`G��"0TX�hQ��q�p8"p��E��8{�ћ]�5¿H.L�[� ߂�պ4p~�0~�11<��>@=`rͳ�6G��M�2#���,ġ�a���f.���9��H�������Y��G��|��%u����q���o��3%7��� ����:*�/L/.��I�J�� 1��73ܸ���	]A�yo�����Ӕ>SO�������޹�����A#-^�+��뺜��|:yݕ`=%��A���/E�8������V�0��A.���lQŇ
B������޲S9���!=X6tB�S ��� ��(��V��`$�ٯ�۲@�w���.�w�K���n��Kv�D�eq�m����-s���9fS?褡����N/#�z�����aS(e��Y�������G+��1�=jeA�䆧��2�.��d�t�d�oI?�fp�d,�|2ߘr!���O�C�5|�c��&p0�g�����ҙ}8DC2�]Ψ�x|��=3Ґ8�+Rn7���U�s��d�|Wa%�۔��C�f�)�=��@��ZUd<��n0t�%���΋�$|ɕ�ɿ*��V󹌷���f��W2�!�3�"�+u%�]�-
�1:'i�a�cF�p�c��)��B�=/<�k���Ʉ ډ�]��p��V��Zl5ZOR��FR��*fOƸ)��SJ]�<��>)��0��^������>'���w�jGp��,�d/�
����r=��?U����"ie��MP�[Tk3G3�e�N��3� V�v�r�ї4h��Sjsº~~�YIB�ˑ-�%|��h-X���b��?|ʎ�yN���n�uX��2٥1�8�%ZG��� ����՘UV�h���,by�+}V�
>��~�1>��v���t+�q�s��(���JySЮ,�+��	ae��8Toe�1���Խ����u���Y�zD��)��^�9̅j����.Di���y�QO�O�7T($���ډ�s��Է����iʠ�);(ۡZ�0��r��YE�������&��#��1������:%��)	�?X��x���X���՞U0�
�/5���C�K���p�� �m���p��ouh�hwϞ�Zc�$��9!"�	) �E�{�I-wi�݀o��
[�]2�X��1%?�1=���vg���Ҵ�<�\wH�9%0
�<s���jfU~��Dnx��)6
w��Ji��^:k�PV	�1�5�7,i�Y�[+`_%q�E�d�_��=���}7
Aڮ��RS�1��Nդ�
X���|�_�*n���'�Zԕ�y�%�WJa<*����QK0��XU㾇0E��k�_�i�i z]!:ZtqΩ5#Бܐ���j�/E��i�HSBf&�UKk�����*|L����6'�ȳ�����{$ɖ�H��Z�T:E�x����M&7��4mG�����5yỉǞ�^x���z}��뺊����2N`��z�d�J���m�	�y������,����/�Mڇ����?%�;k߮	2���{�u/	���	�|��ӴE��u�5��OǄ�r[���Hm z&´nq�Q>��|�4'e�ż��J.������/�.�^j�ǻ%_h���;���`Ł�|�����_�� ��"���w p���}<�C����	�>%qo{�.�30�4����쀇̮�)���I����Cދ)�5�v���W��+��=A�#���������FG8=��V�;�z@%?$�η�}����u���3J��^v�A�`N"�����\1�l�R����=�J'�!~o&�7><܊�n�����Z����y#ڶf�E�{@c�%���D�T�
�q.uْV�w�j�e�j&��p�Q���O$��/������ ��M[L�ZdA�^V��-��nI���ϥ�G8*�ݭ��x�=X�w'_{�HX�~M#_C�'s_�n�H$[ q�E5�^�Ws�:K��$�����v_��B!: ��������{��ꇏH���k�x*��w�c�}rUx���qv-E_`DH@D(DD����)��"riT�ZA�j��웳)���ȶWeA�P�gK.Ȼ�����}�׼���t`���Z'�H#�L�������픑���t�.a����	q�^?I�C8�l/A��Pd��Ϙ1�e�}m�fMՕ"~-��-�~V.��O�x�9�
�	�i�?���=��x�a���!��c]}���V����5�.w��ք��R���q��v�]��> �'G��Z[T������ m=�q�/��=N���y.����"�Ds�Zg��*s����fO����ӷSn.�x�?�|0����)����Ծ�PBe^�V��I+�RXY�M�E����A=bՖu
�#�X��D\"y>�a 9�̿dv�ﾶ����G�?�f���k�ij=�C��fTK@Ԏ�u�n �R)Ԥ5HC��e�*m������'���o (��@�aǚ�d����`/ɪ-Ґ�/�޲Rr���Y���{�[.�g�MD�/��=���LQҢtBؗc=U��	���0\ND���qP���1Ih��Q4Q�K�n�l��N\Rj �

u0�Zi���N{�m7;��v���u�8ܐY�ݠ ϳP��s�(�?b��Gk�0��by瓅��pV�9]LfC�m0@K��]����ZU�FE!��"�A��rz*��"d��i�<W�d�|�nX�#��;�6��"xM	�O���yt=�(� �[9ym�sU���,�v�V��+ƒ�<Y.�_�2�F��|�0/T�Mk[��dns� ���J��7$��-?�]��uy�FT树s09,b���TI�`%��"�	y�\�c/�ǊaD"Xi�ɩ%���9�L�w<#�\�YN,b�(/6����ǃU��R���3�*fd�q��O����0�+��U��:xH�L�|�X�H̠������)�����^P"}�(-���<������͂P�9K��������K�q�����n�Pڈ$�M�����m�t��֮��	S4��,����!�0��b�M�c<AߕH�_���}��޼�Y��#VEk�1�LN����04P_X�
o����B��iX^;K��Z���[����to{�7U5smR��s��q�X���H������#R��)~#Х�\��ǯ�ҟVѭai�;U�����p�P�E��������a�Sg�@��Ws�e���xjm�2M֤̉B������[�=�R�Xvʎ���Gìui�]�pX�p��Z �F���buP�P�����v5&�E��(D@0ꕉ���3�����*��@�!r�yffM�D��g��5�iG]e36���G�6��C����ʚ� >w'�یUv�~N��G{��f62p�J?��~xm���2?;�>|o﷾V�_c�Bs�juek����f�$��M�zkd�_������j��� :�����AW�a����K�uQ�mi�<�O9{�H�|d���|�	(���9�L�)�7��;]�]��K.���@!,z��xP�O�M�;/0m;����
���q_C1�,�y!#D����Ͳ�`g�0ZU��GʐG"�9�8�$�]��:|StFCQ�18�7NlE�,]4�����O��O�Z`�8��u��cm|�0%��'de�1T/��d氡o�g�@�a1k}׶�^��vy.9��&R�|,j�-�e�������N̘��yQ������xC�[��)����+�9�I��p�WH_���Ɓ/SA�@��m���+�S�?����vJX��n��ʶN��^���TJt|��*��K�2��x@; ���m
*�&��T(�g��5�Vvҥ�W�=# �gw�5�H^ -hH�c��C9�I�̴��)���!��u�P9��{1#������(%[�Y%Ǥ�I�1zPG�I�:ȧ*a�Ɗ]�A�+��;�f�}����$�^�zc;�����y-��c�JTo���.ʅx>�� ��w�j.���}�UH���uO�V��}w=rt7}��N}���b� �V��'�p�>������R[���5$ù�X *��Vz}�
H6�1ř��d!��#��ʡe��6��GX�Ezg6H!�h�nc�6�1'���%��h̀��eK|>܃E�}Q^���pl��d���x�x�@R�ݛV�4Ď�U�� ��w6�3�1���R�@Fk���K�S��_4�CS�5�K*�G&A�Q`���ue�m\���wa�[�w��� ֿK�"uw�#�dz�ۢ���B�BWʍ<��r�Qp54�*�H�D�/��P	���]q=`7�fH4tN����X�`���Qt�Kˡ;���uԸ]{��+zp�20S�3�Fj�6�Ķ;F�|ϰEIG�b�iݼ�A0��Y�Jp����C�A,Nk*7D�k}�6�����.ŝ��̛�<IH%r�ꍝ'W��vv%��2>��+�Y;�j��yEڲ%�� �	Q'=t�H�	\�es���qN<�������{.�����(�U'�22݂�q��'�,7���f�Gђ�� %����vըcy/�ܶ��%Ɗ��.���免;�NH�pi�v��γ/vBn�U⡒۟@����{b2�׃�7|����iQ�x���\;��[-��	�wM���c���#��px�u�{� :�����U��&,��}2��ܑ�Z�6x�����M�0x�H�����Q�3>�]��N��4؊
���s}i������lb'm��#r<"��:ۈ�� �'�#����4 ��ǀ��w໧R2+��Ni�@��0S���(¢z#I��T��˨ya�T�(S��OO���Q�O�Ez)������Ǯ��
^`9�����m	rdU�	fT���^��X\Sb��*�`&�'�A��/F�&����0]CF�u���b����`���\(<��jѷ��J҄�Ky������n�Z�uo�7i]����c9z��� L�Q��I�����
�B�V�on��Y��S|��h!ѩ��rk���rd��8X[�$�[�`��',�bҎ\cX���@��$�x�s��k4',j#�'(��:�~�9��ہ�������JD<tj�+�}
�!���8�A�O"���d @��1��rq�Y�qڸA���G�6�ҹ��7��2�$P����9�Hw�-"{��F���7���0�[&�)�9�Y����N]��xE�4s_�tn��!����+�lf+`�s���Ɓ�iÎ,cDI�U���X_th�;�����%�d�r��2�������6Yp��`�����.+_؀*u�A��;��?�H�B��m�i�Ğ�����$/��y��G�R�s_�Q�0O�k/D �������յ#��:�ڰ�v6�p��8a��l���ja��ƕƋxV�U��2L���j���b��� �����%���F�0��X�|+-�N���!n������V������H4IG�cP��ɞ�TvG#�a��Γ~�4]�L$f�V�>N�u?r�1!!Q�f\��j�?$�7�La�I05��Mq�ʓʏ)k��>i�_>�{Z��y9��ܚBZK^e`�����D�S�	:
�4֣���C"����Ŏ`�Y�گnE�I;�nn.��zŭ�
��_���۵����8;�9P�W�{�DD���[iMt��o��G�m��Z�f����p8�� ���n�����]h`$s ��(Ȣa7%
�<�tD �~��c�!-)s}���< ߳�����`�M���@����3����l]={k�Q����K/C}~��[M<x�F��l2g�ڊ���_��6������"��n]�(�"4d+c��!1���ܽ���I��À�6
m�[Au����ې����|!у��K$��w���f~��\��!��Z8������8�v��YW!���:����N('��1qS����SLU6K������U�AY'Q�����j�@E��8����EA��P��S>��D�R%۶{ઞCD
��9�#�x ŋ�~
���J&����r7I!w�H[�M@�8��G@�~�`���90d���QL)�_��׀ðu`�޶�9�A@�M,=��Kq^.u�?Ԁ�r|�lF{�4��nt=�|;F�cـ�#;�`y��l�]�3�_s����ф_�5�WĨ��*�dɖ_s�mǆda4�@��